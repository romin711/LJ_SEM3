<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-97.5525,24.8666,143.953,-94.5048</PageViewport>
<gate>
<ID>2</ID>
<type>AA_AND2</type>
<position>10,-4</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>2,-1</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>2,-7</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>GA_LED</type>
<position>15,-4</position>
<input>
<ID>N_in0</ID>8 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AE_OR2</type>
<position>9,-15.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_TOGGLE</type>
<position>2,-13</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>2,-18</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>-3.5,-3</position>
<gparam>LABEL_TEXT AND</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>-2,-15</position>
<gparam>LABEL_TEXT OR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>GA_LED</type>
<position>15,-15.5</position>
<input>
<ID>N_in0</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AI_XOR2</type>
<position>9,-38</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>1.5,-36</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>1.5,-40</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>30</ID>
<type>GA_LED</type>
<position>14.5,-38</position>
<input>
<ID>N_in0</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>AO_XNOR2</type>
<position>9.5,-49.5</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>34</ID>
<type>BA_NAND2</type>
<position>10.5,5.5</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>36</ID>
<type>BE_NOR2</type>
<position>8.5,-27</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>18 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>37</ID>
<type>AA_LABEL</type>
<position>-4.5,-38</position>
<gparam>LABEL_TEXT X-OR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>38</ID>
<type>AA_TOGGLE</type>
<position>2,-47.5</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>39</ID>
<type>AA_TOGGLE</type>
<position>2,-51.5</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>40</ID>
<type>GA_LED</type>
<position>14.5,-49.5</position>
<input>
<ID>N_in0</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>AA_LABEL</type>
<position>-4.5,-49.5</position>
<gparam>LABEL_TEXT X-NOR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>42</ID>
<type>AA_TOGGLE</type>
<position>2,-24</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_TOGGLE</type>
<position>2,-30</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_LABEL</type>
<position>-3,-26.5</position>
<gparam>LABEL_TEXT NOR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>AA_TOGGLE</type>
<position>2,8</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_TOGGLE</type>
<position>2,3</position>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>47</ID>
<type>AA_LABEL</type>
<position>-2.5,6</position>
<gparam>LABEL_TEXT NAND</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>48</ID>
<type>GA_LED</type>
<position>14.5,-27</position>
<input>
<ID>N_in0</ID>21 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>GA_LED</type>
<position>15,5.5</position>
<input>
<ID>N_in0</ID>22 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5.5,-3,5.5,-1</points>
<intersection>-3 1</intersection>
<intersection>-1 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5.5,-3,7,-3</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>5.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>4,-1,5.5,-1</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>5.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5.5,-7,5.5,-5</points>
<intersection>-7 2</intersection>
<intersection>-5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5.5,-5,7,-5</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>5.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>4,-7,5.5,-7</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>5.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,-14.5,5,-13</points>
<intersection>-14.5 1</intersection>
<intersection>-13 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5,-14.5,6,-14.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>4,-13,5,-13</points>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection>
<intersection>5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,-18,5,-16.5</points>
<intersection>-18 2</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5,-16.5,6,-16.5</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>4,-18,5,-18</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13,-4,14,-4</points>
<connection>
<GID>8</GID>
<name>N_in0</name></connection>
<connection>
<GID>2</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12,-15.5,14,-15.5</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<connection>
<GID>20</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4.5,-37,4.5,-36</points>
<intersection>-37 1</intersection>
<intersection>-36 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4.5,-37,6,-37</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>3.5,-36,4.5,-36</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4.5,-40,4.5,-39</points>
<intersection>-40 2</intersection>
<intersection>-39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4.5,-39,6,-39</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>3.5,-40,4.5,-40</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12,-38,13.5,-38</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<connection>
<GID>30</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,-48.5,5,-47.5</points>
<intersection>-48.5 1</intersection>
<intersection>-47.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5,-48.5,6.5,-48.5</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>4,-47.5,5,-47.5</points>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<intersection>5 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,-51.5,5,-50.5</points>
<intersection>-51.5 2</intersection>
<intersection>-50.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5,-50.5,6.5,-50.5</points>
<connection>
<GID>32</GID>
<name>IN_1</name></connection>
<intersection>5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>4,-51.5,5,-51.5</points>
<connection>
<GID>39</GID>
<name>OUT_0</name></connection>
<intersection>5 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,-49.5,13.5,-49.5</points>
<connection>
<GID>32</GID>
<name>OUT</name></connection>
<connection>
<GID>40</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4.5,-26,4.5,-24</points>
<intersection>-26 1</intersection>
<intersection>-24 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4.5,-26,5.5,-26</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>4,-24,4.5,-24</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4.5,-30,4.5,-28</points>
<intersection>-30 2</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4.5,-28,5.5,-28</points>
<connection>
<GID>36</GID>
<name>IN_1</name></connection>
<intersection>4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>4,-30,4.5,-30</points>
<connection>
<GID>43</GID>
<name>OUT_0</name></connection>
<intersection>4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5.5,6.5,5.5,8</points>
<intersection>6.5 1</intersection>
<intersection>8 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5.5,6.5,7.5,6.5</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>5.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>4,8,5.5,8</points>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection>
<intersection>5.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5.5,3,5.5,4.5</points>
<intersection>3 2</intersection>
<intersection>4.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5.5,4.5,7.5,4.5</points>
<connection>
<GID>34</GID>
<name>IN_1</name></connection>
<intersection>5.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>4,3,5.5,3</points>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection>
<intersection>5.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11.5,-27,13.5,-27</points>
<connection>
<GID>36</GID>
<name>OUT</name></connection>
<connection>
<GID>48</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13.5,5.5,14,5.5</points>
<connection>
<GID>34</GID>
<name>OUT</name></connection>
<connection>
<GID>49</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-4.21111,-10.5111,213.389,-118.067</PageViewport>
<gate>
<ID>51</ID>
<type>AA_LABEL</type>
<position>14.5,-16</position>
<gparam>LABEL_TEXT NAND AS AND</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>BA_NAND2</type>
<position>38,-16.5</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>25 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>54</ID>
<type>BA_NAND2</type>
<position>48.5,-16.5</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>56</ID>
<type>AA_TOGGLE</type>
<position>30,-14</position>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_TOGGLE</type>
<position>30,-19</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>59</ID>
<type>GA_LED</type>
<position>55.5,-16.5</position>
<input>
<ID>N_in0</ID>26 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>14,-37</position>
<gparam>LABEL_TEXT NAND AS OR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>61</ID>
<type>BA_NAND2</type>
<position>38.5,-32.5</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>36 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>62</ID>
<type>BA_NAND2</type>
<position>49,-37.5</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_TOGGLE</type>
<position>29.5,-32.5</position>
<output>
<ID>OUT_0</ID>36 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>65</ID>
<type>GA_LED</type>
<position>56,-37.5</position>
<input>
<ID>N_in0</ID>30 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>BA_NAND2</type>
<position>38.5,-42.5</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>35 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>68</ID>
<type>AA_TOGGLE</type>
<position>29.5,-42.5</position>
<output>
<ID>OUT_0</ID>35 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>69</ID>
<type>AA_LABEL</type>
<position>77.5,-36.5</position>
<gparam>LABEL_TEXT NAND AS NOR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>BA_NAND2</type>
<position>102,-32</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>41 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>71</ID>
<type>BA_NAND2</type>
<position>112.5,-37</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>39 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>72</ID>
<type>AA_TOGGLE</type>
<position>93,-32</position>
<output>
<ID>OUT_0</ID>41 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>74</ID>
<type>BA_NAND2</type>
<position>102,-42</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_1</ID>40 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>75</ID>
<type>AA_TOGGLE</type>
<position>93,-42</position>
<output>
<ID>OUT_0</ID>40 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>76</ID>
<type>BA_NAND2</type>
<position>121.5,-37</position>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>42 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>77</ID>
<type>GA_LED</type>
<position>128.5,-37</position>
<input>
<ID>N_in0</ID>43 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>79</ID>
<type>BA_NAND2</type>
<position>36,-60</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>81</ID>
<type>BA_NAND2</type>
<position>36,-72</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>45 </input>
<output>
<ID>OUT</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>83</ID>
<type>AA_TOGGLE</type>
<position>28.5,-60</position>
<output>
<ID>OUT_0</ID>44 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>84</ID>
<type>AA_TOGGLE</type>
<position>28.5,-72</position>
<output>
<ID>OUT_0</ID>45 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>85</ID>
<type>BA_NAND2</type>
<position>48,-62</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>48 </input>
<output>
<ID>OUT</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>86</ID>
<type>BA_NAND2</type>
<position>48,-70.5</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>45 </input>
<output>
<ID>OUT</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>87</ID>
<type>BA_NAND2</type>
<position>56,-66.5</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>51 </input>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>89</ID>
<type>GA_LED</type>
<position>63,-66.5</position>
<input>
<ID>N_in0</ID>52 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>90</ID>
<type>AA_LABEL</type>
<position>12,-66</position>
<gparam>LABEL_TEXT NAND AS EX-OR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>BA_NAND2</type>
<position>110,-59.5</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>53 </input>
<output>
<ID>OUT</ID>56 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>92</ID>
<type>BA_NAND2</type>
<position>110,-71.5</position>
<input>
<ID>IN_0</ID>54 </input>
<input>
<ID>IN_1</ID>54 </input>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>93</ID>
<type>AA_TOGGLE</type>
<position>102.5,-59.5</position>
<output>
<ID>OUT_0</ID>53 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>94</ID>
<type>AA_TOGGLE</type>
<position>102.5,-71.5</position>
<output>
<ID>OUT_0</ID>54 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>95</ID>
<type>BA_NAND2</type>
<position>122,-61.5</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>55 </input>
<output>
<ID>OUT</ID>57 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>96</ID>
<type>BA_NAND2</type>
<position>122,-70</position>
<input>
<ID>IN_0</ID>56 </input>
<input>
<ID>IN_1</ID>54 </input>
<output>
<ID>OUT</ID>58 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>97</ID>
<type>BA_NAND2</type>
<position>130,-66</position>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>58 </input>
<output>
<ID>OUT</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>99</ID>
<type>AA_LABEL</type>
<position>87.5,-65.5</position>
<gparam>LABEL_TEXT NAND AS EX-NOR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>100</ID>
<type>BA_NAND2</type>
<position>139.5,-66</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>60 </input>
<output>
<ID>OUT</ID>61 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>102</ID>
<type>GA_LED</type>
<position>146.5,-66</position>
<input>
<ID>N_in0</ID>61 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,-17.5,45.5,-15.5</points>
<connection>
<GID>54</GID>
<name>IN_1</name></connection>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-16.5,45.5,-16.5</points>
<connection>
<GID>53</GID>
<name>OUT</name></connection>
<intersection>45.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-15.5,33.5,-14</points>
<intersection>-15.5 1</intersection>
<intersection>-14 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-15.5,35,-15.5</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>33.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,-14,33.5,-14</points>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection>
<intersection>33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-19,33.5,-17.5</points>
<intersection>-19 2</intersection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-17.5,35,-17.5</points>
<connection>
<GID>53</GID>
<name>IN_1</name></connection>
<intersection>33.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,-19,33.5,-19</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<intersection>33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>51.5,-16.5,54.5,-16.5</points>
<connection>
<GID>59</GID>
<name>N_in0</name></connection>
<connection>
<GID>54</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>52,-37.5,55,-37.5</points>
<connection>
<GID>62</GID>
<name>OUT</name></connection>
<connection>
<GID>65</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-36.5,43.5,-32.5</points>
<intersection>-36.5 1</intersection>
<intersection>-32.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-36.5,46,-36.5</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>43.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>41.5,-32.5,43.5,-32.5</points>
<connection>
<GID>61</GID>
<name>OUT</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-42.5,43.5,-38.5</points>
<intersection>-42.5 2</intersection>
<intersection>-38.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-38.5,46,-38.5</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<intersection>43.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>41.5,-42.5,43.5,-42.5</points>
<connection>
<GID>66</GID>
<name>OUT</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-43.5,35.5,-41.5</points>
<connection>
<GID>66</GID>
<name>IN_1</name></connection>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>-42.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-42.5,35.5,-42.5</points>
<connection>
<GID>68</GID>
<name>OUT_0</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-33.5,35.5,-31.5</points>
<connection>
<GID>61</GID>
<name>IN_1</name></connection>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-32.5,35.5,-32.5</points>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-36,107,-32</points>
<intersection>-36 1</intersection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-36,109.5,-36</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<intersection>107 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>105,-32,107,-32</points>
<connection>
<GID>70</GID>
<name>OUT</name></connection>
<intersection>107 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-42,107,-38</points>
<intersection>-42 2</intersection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-38,109.5,-38</points>
<connection>
<GID>71</GID>
<name>IN_1</name></connection>
<intersection>107 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>105,-42,107,-42</points>
<connection>
<GID>74</GID>
<name>OUT</name></connection>
<intersection>107 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-43,99,-41</points>
<connection>
<GID>74</GID>
<name>IN_1</name></connection>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>-42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95,-42,99,-42</points>
<connection>
<GID>75</GID>
<name>OUT_0</name></connection>
<intersection>99 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-33,99,-31</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95,-32,99,-32</points>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection>
<intersection>99 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118.5,-38,118.5,-36</points>
<connection>
<GID>76</GID>
<name>IN_1</name></connection>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>-37 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>115.5,-37,118.5,-37</points>
<connection>
<GID>71</GID>
<name>OUT</name></connection>
<intersection>118.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124.5,-37,127.5,-37</points>
<connection>
<GID>76</GID>
<name>OUT</name></connection>
<connection>
<GID>77</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-61,33,-55.5</points>
<connection>
<GID>79</GID>
<name>IN_1</name></connection>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>-60 1</intersection>
<intersection>-55.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-60,33,-60</points>
<connection>
<GID>83</GID>
<name>OUT_0</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33,-55.5,45,-55.5</points>
<intersection>33 0</intersection>
<intersection>45 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>45,-61,45,-55.5</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<intersection>-55.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-76.5,33,-71</points>
<connection>
<GID>81</GID>
<name>IN_1</name></connection>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<intersection>-76.5 2</intersection>
<intersection>-72 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-72,33,-72</points>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33,-76.5,45,-76.5</points>
<intersection>33 0</intersection>
<intersection>45 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>45,-76.5,45,-71.5</points>
<connection>
<GID>86</GID>
<name>IN_1</name></connection>
<intersection>-76.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-72,42.5,-63</points>
<intersection>-72 2</intersection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42.5,-63,45,-63</points>
<connection>
<GID>85</GID>
<name>IN_1</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>39,-72,42.5,-72</points>
<connection>
<GID>81</GID>
<name>OUT</name></connection>
<intersection>42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,-69.5,42,-60</points>
<intersection>-69.5 1</intersection>
<intersection>-60 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42,-69.5,45,-69.5</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<intersection>42 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>39,-60,42,-60</points>
<connection>
<GID>79</GID>
<name>OUT</name></connection>
<intersection>42 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-65.5,52,-62</points>
<intersection>-65.5 1</intersection>
<intersection>-62 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52,-65.5,53,-65.5</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51,-62,52,-62</points>
<connection>
<GID>85</GID>
<name>OUT</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-70.5,52,-67.5</points>
<intersection>-70.5 2</intersection>
<intersection>-67.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52,-67.5,53,-67.5</points>
<connection>
<GID>87</GID>
<name>IN_1</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51,-70.5,52,-70.5</points>
<connection>
<GID>86</GID>
<name>OUT</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59,-66.5,62,-66.5</points>
<connection>
<GID>87</GID>
<name>OUT</name></connection>
<connection>
<GID>89</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-60.5,107,-54.5</points>
<connection>
<GID>91</GID>
<name>IN_1</name></connection>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>-59.5 1</intersection>
<intersection>-54.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,-59.5,107,-59.5</points>
<connection>
<GID>93</GID>
<name>OUT_0</name></connection>
<intersection>107 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>107,-54.5,119,-54.5</points>
<intersection>107 0</intersection>
<intersection>119 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>119,-60.5,119,-54.5</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<intersection>-54.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-76,107,-70.5</points>
<connection>
<GID>92</GID>
<name>IN_1</name></connection>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<intersection>-76 2</intersection>
<intersection>-71.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104.5,-71.5,107,-71.5</points>
<connection>
<GID>94</GID>
<name>OUT_0</name></connection>
<intersection>107 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>107,-76,119,-76</points>
<intersection>107 0</intersection>
<intersection>119 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>119,-76,119,-71</points>
<connection>
<GID>96</GID>
<name>IN_1</name></connection>
<intersection>-76 2</intersection></vsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117,-71.5,117,-62.5</points>
<intersection>-71.5 3</intersection>
<intersection>-62.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117,-62.5,119,-62.5</points>
<connection>
<GID>95</GID>
<name>IN_1</name></connection>
<intersection>117 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>113,-71.5,117,-71.5</points>
<connection>
<GID>92</GID>
<name>OUT</name></connection>
<intersection>117 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116,-69,116,-59.5</points>
<intersection>-69 1</intersection>
<intersection>-59.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116,-69,119,-69</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>116 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113,-59.5,116,-59.5</points>
<connection>
<GID>91</GID>
<name>OUT</name></connection>
<intersection>116 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126,-65,126,-61.5</points>
<intersection>-65 1</intersection>
<intersection>-61.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126,-65,127,-65</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>126 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>125,-61.5,126,-61.5</points>
<connection>
<GID>95</GID>
<name>OUT</name></connection>
<intersection>126 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126,-70,126,-67</points>
<intersection>-70 2</intersection>
<intersection>-67 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126,-67,127,-67</points>
<connection>
<GID>97</GID>
<name>IN_1</name></connection>
<intersection>126 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>125,-70,126,-70</points>
<connection>
<GID>96</GID>
<name>OUT</name></connection>
<intersection>126 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136.5,-67,136.5,-65</points>
<connection>
<GID>100</GID>
<name>IN_1</name></connection>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>-66 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133,-66,136.5,-66</points>
<connection>
<GID>97</GID>
<name>OUT</name></connection>
<intersection>136.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142.5,-66,145.5,-66</points>
<connection>
<GID>102</GID>
<name>N_in0</name></connection>
<connection>
<GID>100</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>-24.3491,11.7502,166.551,-82.608</PageViewport>
<gate>
<ID>104</ID>
<type>BE_NOR2</type>
<position>31,-11</position>
<input>
<ID>IN_0</ID>62 </input>
<input>
<ID>IN_1</ID>62 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>106</ID>
<type>AA_TOGGLE</type>
<position>24,-11</position>
<output>
<ID>OUT_0</ID>62 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>108</ID>
<type>GA_LED</type>
<position>36.5,-11</position>
<input>
<ID>N_in0</ID>63 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>110</ID>
<type>AA_LABEL</type>
<position>12.5,-10.5</position>
<gparam>LABEL_TEXT NOR AS NOT</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>111</ID>
<type>BE_NOR2</type>
<position>27,-24.5</position>
<input>
<ID>IN_0</ID>74 </input>
<input>
<ID>IN_1</ID>75 </input>
<output>
<ID>OUT</ID>73 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>112</ID>
<type>BE_NOR2</type>
<position>33.5,-24.5</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>73 </input>
<output>
<ID>OUT</ID>76 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>113</ID>
<type>BE_NOR2</type>
<position>31,-46.5</position>
<input>
<ID>IN_0</ID>78 </input>
<input>
<ID>IN_1</ID>78 </input>
<output>
<ID>OUT</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>114</ID>
<type>BE_NOR2</type>
<position>31,-36</position>
<input>
<ID>IN_0</ID>77 </input>
<input>
<ID>IN_1</ID>77 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>115</ID>
<type>BE_NOR2</type>
<position>106,-11.5</position>
<input>
<ID>IN_0</ID>89 </input>
<input>
<ID>IN_1</ID>89 </input>
<output>
<ID>OUT</ID>94 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>116</ID>
<type>BE_NOR2</type>
<position>42,-41.5</position>
<input>
<ID>IN_0</ID>80 </input>
<input>
<ID>IN_1</ID>79 </input>
<output>
<ID>OUT</ID>81 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>118</ID>
<type>BE_NOR2</type>
<position>106.5,-22</position>
<input>
<ID>IN_0</ID>90 </input>
<input>
<ID>IN_1</ID>90 </input>
<output>
<ID>OUT</ID>93 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>119</ID>
<type>GA_LED</type>
<position>38.5,-24.5</position>
<input>
<ID>N_in0</ID>76 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>120</ID>
<type>AA_TOGGLE</type>
<position>19,-22.5</position>
<output>
<ID>OUT_0</ID>74 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>121</ID>
<type>AA_TOGGLE</type>
<position>19,-27</position>
<output>
<ID>OUT_0</ID>75 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>122</ID>
<type>AA_LABEL</type>
<position>7.5,-24.5</position>
<gparam>LABEL_TEXT NOR AS OR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>124</ID>
<type>AA_TOGGLE</type>
<position>19.5,-36</position>
<output>
<ID>OUT_0</ID>77 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>126</ID>
<type>AA_TOGGLE</type>
<position>19.5,-46.5</position>
<output>
<ID>OUT_0</ID>78 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>128</ID>
<type>GA_LED</type>
<position>48.5,-41.5</position>
<input>
<ID>N_in0</ID>81 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>131</ID>
<type>AA_LABEL</type>
<position>8.5,-41</position>
<gparam>LABEL_TEXT NOR AS AND</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>132</ID>
<type>BE_NOR2</type>
<position>31.5,-68</position>
<input>
<ID>IN_0</ID>83 </input>
<input>
<ID>IN_1</ID>83 </input>
<output>
<ID>OUT</ID>84 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>133</ID>
<type>BE_NOR2</type>
<position>31.5,-57.5</position>
<input>
<ID>IN_0</ID>82 </input>
<input>
<ID>IN_1</ID>82 </input>
<output>
<ID>OUT</ID>85 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>134</ID>
<type>BE_NOR2</type>
<position>42.5,-63</position>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>84 </input>
<output>
<ID>OUT</ID>87 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>135</ID>
<type>AA_TOGGLE</type>
<position>20,-57.5</position>
<output>
<ID>OUT_0</ID>82 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>136</ID>
<type>AA_TOGGLE</type>
<position>20,-68</position>
<output>
<ID>OUT_0</ID>83 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>138</ID>
<type>AA_LABEL</type>
<position>9,-63</position>
<gparam>LABEL_TEXT NOR AS NAND</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>139</ID>
<type>BE_NOR2</type>
<position>51.5,-63</position>
<input>
<ID>IN_0</ID>87 </input>
<input>
<ID>IN_1</ID>87 </input>
<output>
<ID>OUT</ID>88 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>140</ID>
<type>GA_LED</type>
<position>57.5,-63</position>
<input>
<ID>N_in0</ID>88 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>142</ID>
<type>AA_TOGGLE</type>
<position>97,-11.5</position>
<output>
<ID>OUT_0</ID>89 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>143</ID>
<type>AA_TOGGLE</type>
<position>97.5,-22</position>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>145</ID>
<type>BE_NOR2</type>
<position>118.5,-13.5</position>
<input>
<ID>IN_0</ID>89 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>95 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>146</ID>
<type>BE_NOR2</type>
<position>119,-20.5</position>
<input>
<ID>IN_0</ID>94 </input>
<input>
<ID>IN_1</ID>90 </input>
<output>
<ID>OUT</ID>96 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>147</ID>
<type>BE_NOR2</type>
<position>127.5,-17</position>
<input>
<ID>IN_0</ID>95 </input>
<input>
<ID>IN_1</ID>96 </input>
<output>
<ID>OUT</ID>108 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>150</ID>
<type>AA_LABEL</type>
<position>91.5,-16.5</position>
<gparam>LABEL_TEXT NOR AS X-OR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>151</ID>
<type>BE_NOR2</type>
<position>105.5,-43.5</position>
<input>
<ID>IN_0</ID>112 </input>
<input>
<ID>IN_1</ID>112 </input>
<output>
<ID>OUT</ID>110 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>152</ID>
<type>BE_NOR2</type>
<position>106,-54</position>
<input>
<ID>IN_0</ID>113 </input>
<input>
<ID>IN_1</ID>113 </input>
<output>
<ID>OUT</ID>111 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>153</ID>
<type>AA_TOGGLE</type>
<position>96.5,-43.5</position>
<output>
<ID>OUT_0</ID>112 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>154</ID>
<type>AA_TOGGLE</type>
<position>96.5,-54</position>
<output>
<ID>OUT_0</ID>113 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>155</ID>
<type>BE_NOR2</type>
<position>118,-45.5</position>
<input>
<ID>IN_0</ID>110 </input>
<input>
<ID>IN_1</ID>111 </input>
<output>
<ID>OUT</ID>102 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>156</ID>
<type>BE_NOR2</type>
<position>118.5,-52.5</position>
<input>
<ID>IN_0</ID>112 </input>
<input>
<ID>IN_1</ID>113 </input>
<output>
<ID>OUT</ID>103 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>157</ID>
<type>BE_NOR2</type>
<position>127,-49</position>
<input>
<ID>IN_0</ID>102 </input>
<input>
<ID>IN_1</ID>103 </input>
<output>
<ID>OUT</ID>105 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>159</ID>
<type>AA_LABEL</type>
<position>88.5,-49</position>
<gparam>LABEL_TEXT NOR AS X-NOR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>160</ID>
<type>BE_NOR2</type>
<position>134.5,-49</position>
<input>
<ID>IN_0</ID>105 </input>
<input>
<ID>IN_1</ID>105 </input>
<output>
<ID>OUT</ID>107 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>165</ID>
<type>GA_LED</type>
<position>140,-49</position>
<input>
<ID>N_in0</ID>107 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>166</ID>
<type>BE_NOR2</type>
<position>136.5,-17</position>
<input>
<ID>IN_0</ID>108 </input>
<input>
<ID>IN_1</ID>108 </input>
<output>
<ID>OUT</ID>109 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>168</ID>
<type>GA_LED</type>
<position>142,-17</position>
<input>
<ID>N_in0</ID>109 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-12,28,-10</points>
<connection>
<GID>104</GID>
<name>IN_1</name></connection>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-11,28,-11</points>
<connection>
<GID>106</GID>
<name>OUT_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-11,35.5,-11</points>
<connection>
<GID>108</GID>
<name>N_in0</name></connection>
<connection>
<GID>104</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-25.5,30.5,-23.5</points>
<connection>
<GID>112</GID>
<name>IN_1</name></connection>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-24.5,30.5,-24.5</points>
<connection>
<GID>111</GID>
<name>OUT</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-23.5,22.5,-22.5</points>
<intersection>-23.5 1</intersection>
<intersection>-22.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-23.5,24,-23.5</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21,-22.5,22.5,-22.5</points>
<connection>
<GID>120</GID>
<name>OUT_0</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-27,22.5,-25.5</points>
<intersection>-27 2</intersection>
<intersection>-25.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-25.5,24,-25.5</points>
<connection>
<GID>111</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21,-27,22.5,-27</points>
<connection>
<GID>121</GID>
<name>OUT_0</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36.5,-24.5,37.5,-24.5</points>
<connection>
<GID>112</GID>
<name>OUT</name></connection>
<connection>
<GID>119</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-37,28,-35</points>
<connection>
<GID>114</GID>
<name>IN_1</name></connection>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21.5,-36,28,-36</points>
<connection>
<GID>124</GID>
<name>OUT_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-47.5,28,-45.5</points>
<connection>
<GID>113</GID>
<name>IN_1</name></connection>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>-46.5 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>21.5,-46.5,28,-46.5</points>
<connection>
<GID>126</GID>
<name>OUT_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-46.5,36.5,-42.5</points>
<intersection>-46.5 2</intersection>
<intersection>-42.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36.5,-42.5,39,-42.5</points>
<connection>
<GID>116</GID>
<name>IN_1</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-46.5,36.5,-46.5</points>
<connection>
<GID>113</GID>
<name>OUT</name></connection>
<intersection>36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-40.5,36.5,-36</points>
<intersection>-40.5 1</intersection>
<intersection>-36 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36.5,-40.5,39,-40.5</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-36,36.5,-36</points>
<connection>
<GID>114</GID>
<name>OUT</name></connection>
<intersection>36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-41.5,47.5,-41.5</points>
<connection>
<GID>128</GID>
<name>N_in0</name></connection>
<intersection>45 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>45,-41.5,45,-41.5</points>
<connection>
<GID>116</GID>
<name>OUT</name></connection>
<intersection>-41.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-58.5,28.5,-56.5</points>
<connection>
<GID>133</GID>
<name>IN_1</name></connection>
<connection>
<GID>133</GID>
<name>IN_0</name></connection>
<intersection>-57.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-57.5,28.5,-57.5</points>
<connection>
<GID>135</GID>
<name>OUT_0</name></connection>
<intersection>28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-69,28.5,-67</points>
<connection>
<GID>132</GID>
<name>IN_1</name></connection>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>-68 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>22,-68,28.5,-68</points>
<connection>
<GID>136</GID>
<name>OUT_0</name></connection>
<intersection>28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-68,37,-64</points>
<intersection>-68 2</intersection>
<intersection>-64 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-64,39.5,-64</points>
<connection>
<GID>134</GID>
<name>IN_1</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-68,37,-68</points>
<connection>
<GID>132</GID>
<name>OUT</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-62,37,-57.5</points>
<intersection>-62 1</intersection>
<intersection>-57.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-62,39.5,-62</points>
<connection>
<GID>134</GID>
<name>IN_0</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-57.5,37,-57.5</points>
<connection>
<GID>133</GID>
<name>OUT</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48.5,-64,48.5,-62</points>
<connection>
<GID>139</GID>
<name>IN_1</name></connection>
<connection>
<GID>139</GID>
<name>IN_0</name></connection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45.5,-63,48.5,-63</points>
<connection>
<GID>134</GID>
<name>OUT</name></connection>
<intersection>48.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54.5,-63,56.5,-63</points>
<connection>
<GID>139</GID>
<name>OUT</name></connection>
<connection>
<GID>140</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103,-12.5,103,-6.5</points>
<connection>
<GID>115</GID>
<name>IN_1</name></connection>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<intersection>-11.5 1</intersection>
<intersection>-6.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99,-11.5,103,-11.5</points>
<connection>
<GID>142</GID>
<name>OUT_0</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-6.5,115.5,-6.5</points>
<intersection>103 0</intersection>
<intersection>115.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>115.5,-12.5,115.5,-6.5</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<intersection>-6.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103.5,-27,103.5,-21</points>
<connection>
<GID>118</GID>
<name>IN_1</name></connection>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>-27 2</intersection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99.5,-22,103.5,-22</points>
<connection>
<GID>143</GID>
<name>OUT_0</name></connection>
<intersection>103.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,-27,116,-27</points>
<intersection>103.5 0</intersection>
<intersection>116 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>116,-27,116,-21.5</points>
<connection>
<GID>146</GID>
<name>IN_1</name></connection>
<intersection>-27 2</intersection></vsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-22,111,-14.5</points>
<intersection>-22 2</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111,-14.5,115.5,-14.5</points>
<connection>
<GID>145</GID>
<name>IN_1</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>109.5,-22,111,-22</points>
<connection>
<GID>118</GID>
<name>OUT</name></connection>
<intersection>111 0</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112.5,-19.5,112.5,-11.5</points>
<intersection>-19.5 1</intersection>
<intersection>-11.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112.5,-19.5,116,-19.5</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<intersection>112.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>109,-11.5,112.5,-11.5</points>
<connection>
<GID>115</GID>
<name>OUT</name></connection>
<intersection>112.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123,-16,123,-13.5</points>
<intersection>-16 1</intersection>
<intersection>-13.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123,-16,124.5,-16</points>
<connection>
<GID>147</GID>
<name>IN_0</name></connection>
<intersection>123 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>121.5,-13.5,123,-13.5</points>
<connection>
<GID>145</GID>
<name>OUT</name></connection>
<intersection>123 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123,-20.5,123,-18</points>
<intersection>-20.5 2</intersection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123,-18,124.5,-18</points>
<connection>
<GID>147</GID>
<name>IN_1</name></connection>
<intersection>123 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>122,-20.5,123,-20.5</points>
<connection>
<GID>146</GID>
<name>OUT</name></connection>
<intersection>123 0</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,-48,122.5,-45.5</points>
<intersection>-48 1</intersection>
<intersection>-45.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122.5,-48,124,-48</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>122.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>121,-45.5,122.5,-45.5</points>
<connection>
<GID>155</GID>
<name>OUT</name></connection>
<intersection>122.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,-52.5,122.5,-50</points>
<intersection>-52.5 2</intersection>
<intersection>-50 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122.5,-50,124,-50</points>
<connection>
<GID>157</GID>
<name>IN_1</name></connection>
<intersection>122.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>121.5,-52.5,122.5,-52.5</points>
<connection>
<GID>156</GID>
<name>OUT</name></connection>
<intersection>122.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131.5,-50,131.5,-48</points>
<connection>
<GID>160</GID>
<name>IN_1</name></connection>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<intersection>-49 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130,-49,131.5,-49</points>
<connection>
<GID>157</GID>
<name>OUT</name></connection>
<intersection>131.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>137.5,-49,139,-49</points>
<connection>
<GID>160</GID>
<name>OUT</name></connection>
<connection>
<GID>165</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133.5,-18,133.5,-16</points>
<connection>
<GID>166</GID>
<name>IN_1</name></connection>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130.5,-17,133.5,-17</points>
<connection>
<GID>147</GID>
<name>OUT</name></connection>
<intersection>133.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>139.5,-17,141,-17</points>
<connection>
<GID>168</GID>
<name>N_in0</name></connection>
<connection>
<GID>166</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111.5,-44.5,111.5,-43.5</points>
<intersection>-44.5 1</intersection>
<intersection>-43.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111.5,-44.5,115,-44.5</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<intersection>111.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>108.5,-43.5,111.5,-43.5</points>
<connection>
<GID>151</GID>
<name>OUT</name></connection>
<intersection>111.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,-54,112,-46.5</points>
<intersection>-54 2</intersection>
<intersection>-46.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112,-46.5,115,-46.5</points>
<connection>
<GID>155</GID>
<name>IN_1</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>109,-54,112,-54</points>
<connection>
<GID>152</GID>
<name>OUT</name></connection>
<intersection>112 0</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102.5,-49,102.5,-42.5</points>
<connection>
<GID>151</GID>
<name>IN_1</name></connection>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<intersection>-49 2</intersection>
<intersection>-43.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98.5,-43.5,102.5,-43.5</points>
<connection>
<GID>153</GID>
<name>OUT_0</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>102.5,-49,115.5,-49</points>
<intersection>102.5 0</intersection>
<intersection>115.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>115.5,-51.5,115.5,-49</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<intersection>-49 2</intersection></vsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103,-59,103,-53</points>
<connection>
<GID>152</GID>
<name>IN_1</name></connection>
<connection>
<GID>152</GID>
<name>IN_0</name></connection>
<intersection>-59 2</intersection>
<intersection>-54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98.5,-54,103,-54</points>
<connection>
<GID>154</GID>
<name>OUT_0</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103,-59,115.5,-59</points>
<intersection>103 0</intersection>
<intersection>115.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>115.5,-59,115.5,-53.5</points>
<connection>
<GID>156</GID>
<name>IN_1</name></connection>
<intersection>-59 2</intersection></vsegment></shape></wire></page 2>
<page 3>
<PageViewport>-220.805,29.5697,208.538,-182.646</PageViewport>
<gate>
<ID>193</ID>
<type>GA_LED</type>
<position>14,-24.5</position>
<input>
<ID>N_in0</ID>123 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>195</ID>
<type>AA_INVERTER</type>
<position>67.5,-1</position>
<input>
<ID>IN_0</ID>128 </input>
<output>
<ID>OUT_0</ID>130 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>197</ID>
<type>AA_INVERTER</type>
<position>69,-17.5</position>
<input>
<ID>IN_0</ID>129 </input>
<output>
<ID>OUT_0</ID>131 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>198</ID>
<type>AA_LABEL</type>
<position>58,-1</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>199</ID>
<type>AA_LABEL</type>
<position>58.5,-17</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>201</ID>
<type>AA_TOGGLE</type>
<position>61,-1</position>
<output>
<ID>OUT_0</ID>128 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>202</ID>
<type>AA_TOGGLE</type>
<position>61.5,-17.5</position>
<output>
<ID>OUT_0</ID>129 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>204</ID>
<type>AA_AND2</type>
<position>82,2.5</position>
<input>
<ID>IN_0</ID>130 </input>
<input>
<ID>IN_1</ID>129 </input>
<output>
<ID>OUT</ID>134 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>206</ID>
<type>AA_AND2</type>
<position>82.5,-10</position>
<input>
<ID>IN_0</ID>128 </input>
<input>
<ID>IN_1</ID>131 </input>
<output>
<ID>OUT</ID>133 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>208</ID>
<type>AA_AND2</type>
<position>83,-24</position>
<input>
<ID>IN_0</ID>128 </input>
<input>
<ID>IN_1</ID>129 </input>
<output>
<ID>OUT</ID>132 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>210</ID>
<type>AE_OR2</type>
<position>91.5,-4.5</position>
<input>
<ID>IN_0</ID>134 </input>
<input>
<ID>IN_1</ID>133 </input>
<output>
<ID>OUT</ID>135 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>212</ID>
<type>GA_LED</type>
<position>88.5,-24</position>
<input>
<ID>N_in0</ID>132 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>214</ID>
<type>GA_LED</type>
<position>96.5,-4.5</position>
<input>
<ID>N_in0</ID>135 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>215</ID>
<type>AA_LABEL</type>
<position>72,12.5</position>
<gparam>LABEL_TEXT HALF ADDER USING AOI</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>217</ID>
<type>AA_LABEL</type>
<position>22.5,-10</position>
<gparam>LABEL_TEXT CARRY</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>218</ID>
<type>AA_LABEL</type>
<position>23.5,-25</position>
<gparam>LABEL_TEXT SUM</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>219</ID>
<type>AA_LABEL</type>
<position>104.5,-4.5</position>
<gparam>LABEL_TEXT CARRY</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>220</ID>
<type>AA_LABEL</type>
<position>93.5,-23.5</position>
<gparam>LABEL_TEXT SUM</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>221</ID>
<type>AA_LABEL</type>
<position>-15.5,-54.5</position>
<gparam>LABEL_TEXT HALF ADDER USING NOR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>223</ID>
<type>BE_NOR2</type>
<position>-30.5,-70.5</position>
<input>
<ID>IN_0</ID>136 </input>
<input>
<ID>IN_1</ID>136 </input>
<output>
<ID>OUT</ID>139 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>224</ID>
<type>BE_NOR2</type>
<position>-30.5,-86</position>
<input>
<ID>IN_0</ID>137 </input>
<input>
<ID>IN_1</ID>137 </input>
<output>
<ID>OUT</ID>138 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>225</ID>
<type>BE_NOR2</type>
<position>-14.5,-65.5</position>
<input>
<ID>IN_0</ID>136 </input>
<input>
<ID>IN_1</ID>138 </input>
<output>
<ID>OUT</ID>140 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>226</ID>
<type>BE_NOR2</type>
<position>-14,-78.5</position>
<input>
<ID>IN_0</ID>139 </input>
<input>
<ID>IN_1</ID>137 </input>
<output>
<ID>OUT</ID>141 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>227</ID>
<type>BE_NOR2</type>
<position>-14,-92</position>
<input>
<ID>IN_0</ID>139 </input>
<input>
<ID>IN_1</ID>138 </input>
<output>
<ID>OUT</ID>142 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>228</ID>
<type>BE_NOR2</type>
<position>4.5,-72</position>
<input>
<ID>IN_0</ID>140 </input>
<input>
<ID>IN_1</ID>141 </input>
<output>
<ID>OUT</ID>143 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>233</ID>
<type>AA_TOGGLE</type>
<position>-37.5,-70.5</position>
<output>
<ID>OUT_0</ID>136 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>234</ID>
<type>AA_TOGGLE</type>
<position>-37,-86</position>
<output>
<ID>OUT_0</ID>137 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>236</ID>
<type>GA_LED</type>
<position>-9,-92</position>
<input>
<ID>N_in0</ID>142 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>238</ID>
<type>GA_LED</type>
<position>9.5,-72</position>
<input>
<ID>N_in0</ID>143 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>170</ID>
<type>BA_NAND2</type>
<position>-30.5,-8.5</position>
<input>
<ID>IN_0</ID>124 </input>
<input>
<ID>IN_1</ID>124 </input>
<output>
<ID>OUT</ID>126 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>171</ID>
<type>BA_NAND2</type>
<position>-30.5,-24</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>125 </input>
<output>
<ID>OUT</ID>127 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>173</ID>
<type>AA_LABEL</type>
<position>-22.5,13.5</position>
<gparam>LABEL_TEXT HALF ADDER USING NAND</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>175</ID>
<type>BA_NAND2</type>
<position>-11.5,-3.5</position>
<input>
<ID>IN_0</ID>124 </input>
<input>
<ID>IN_1</ID>125 </input>
<output>
<ID>OUT</ID>121 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>177</ID>
<type>BA_NAND2</type>
<position>-11.5,-17.5</position>
<input>
<ID>IN_0</ID>126 </input>
<input>
<ID>IN_1</ID>125 </input>
<output>
<ID>OUT</ID>119 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>178</ID>
<type>BA_NAND2</type>
<position>-11.5,-30.5</position>
<input>
<ID>IN_0</ID>124 </input>
<input>
<ID>IN_1</ID>127 </input>
<output>
<ID>OUT</ID>120 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>180</ID>
<type>BA_NAND2</type>
<position>8,-9.5</position>
<input>
<ID>IN_0</ID>121 </input>
<input>
<ID>IN_1</ID>121 </input>
<output>
<ID>OUT</ID>122 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>181</ID>
<type>BA_NAND2</type>
<position>9,-24.5</position>
<input>
<ID>IN_0</ID>119 </input>
<input>
<ID>IN_1</ID>120 </input>
<output>
<ID>OUT</ID>123 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>183</ID>
<type>AA_TOGGLE</type>
<position>-42.5,-8.5</position>
<output>
<ID>OUT_0</ID>124 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>185</ID>
<type>AA_TOGGLE</type>
<position>-42,-24</position>
<output>
<ID>OUT_0</ID>125 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>187</ID>
<type>AA_LABEL</type>
<position>-46.5,-8</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>188</ID>
<type>AA_LABEL</type>
<position>-45.5,-23.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>192</ID>
<type>GA_LED</type>
<position>13,-9.5</position>
<input>
<ID>N_in0</ID>122 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1.5,-23.5,-1.5,-17.5</points>
<intersection>-23.5 1</intersection>
<intersection>-17.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1.5,-23.5,6,-23.5</points>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<intersection>-1.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-8.5,-17.5,-1.5,-17.5</points>
<connection>
<GID>177</GID>
<name>OUT</name></connection>
<intersection>-1.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1.5,-30.5,-1.5,-25.5</points>
<intersection>-30.5 2</intersection>
<intersection>-25.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1.5,-25.5,6,-25.5</points>
<connection>
<GID>181</GID>
<name>IN_1</name></connection>
<intersection>-1.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-8.5,-30.5,-1.5,-30.5</points>
<connection>
<GID>178</GID>
<name>OUT</name></connection>
<intersection>-1.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,-10.5,5,-8.5</points>
<connection>
<GID>180</GID>
<name>IN_1</name></connection>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<intersection>-9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-8.5,-9.5,5,-9.5</points>
<intersection>-8.5 2</intersection>
<intersection>5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-8.5,-9.5,-8.5,-3.5</points>
<connection>
<GID>175</GID>
<name>OUT</name></connection>
<intersection>-9.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11,-9.5,12,-9.5</points>
<connection>
<GID>180</GID>
<name>OUT</name></connection>
<connection>
<GID>192</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12,-24.5,13,-24.5</points>
<connection>
<GID>193</GID>
<name>N_in0</name></connection>
<connection>
<GID>181</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33.5,-9.5,-33.5,-2.5</points>
<connection>
<GID>170</GID>
<name>IN_1</name></connection>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>-8.5 1</intersection>
<intersection>-2.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-40.5,-8.5,-33.5,-8.5</points>
<connection>
<GID>183</GID>
<name>OUT_0</name></connection>
<intersection>-33.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-33.5,-2.5,-14.5,-2.5</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>-33.5 0</intersection>
<intersection>-18 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-18,-29.5,-18,-2.5</points>
<intersection>-29.5 4</intersection>
<intersection>-2.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-18,-29.5,-14.5,-29.5</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<intersection>-18 3</intersection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36,-25,-36,-4.5</points>
<intersection>-25 3</intersection>
<intersection>-24 1</intersection>
<intersection>-23 4</intersection>
<intersection>-4.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-40,-24,-36,-24</points>
<connection>
<GID>185</GID>
<name>OUT_0</name></connection>
<intersection>-36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-36,-4.5,-14.5,-4.5</points>
<connection>
<GID>175</GID>
<name>IN_1</name></connection>
<intersection>-36 0</intersection>
<intersection>-25.5 5</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-36,-25,-33.5,-25</points>
<connection>
<GID>171</GID>
<name>IN_1</name></connection>
<intersection>-36 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-36,-23,-33.5,-23</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<intersection>-36 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-25.5,-18.5,-25.5,-4.5</points>
<intersection>-18.5 6</intersection>
<intersection>-4.5 2</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-25.5,-18.5,-14.5,-18.5</points>
<connection>
<GID>177</GID>
<name>IN_1</name></connection>
<intersection>-25.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-21,-16.5,-21,-8.5</points>
<intersection>-16.5 1</intersection>
<intersection>-8.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-21,-16.5,-14.5,-16.5</points>
<connection>
<GID>177</GID>
<name>IN_0</name></connection>
<intersection>-21 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-27.5,-8.5,-21,-8.5</points>
<connection>
<GID>170</GID>
<name>OUT</name></connection>
<intersection>-21 0</intersection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-21,-31.5,-21,-24</points>
<intersection>-31.5 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-27.5,-24,-21,-24</points>
<connection>
<GID>171</GID>
<name>OUT</name></connection>
<intersection>-21 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-31.5,-14.5,-31.5</points>
<connection>
<GID>178</GID>
<name>IN_1</name></connection>
<intersection>-21 0</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>63,-5.5,76.5,-5.5</points>
<intersection>63 4</intersection>
<intersection>64.5 3</intersection>
<intersection>76.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>76.5,-23,76.5,-5.5</points>
<intersection>-23 6</intersection>
<intersection>-9 12</intersection>
<intersection>-5.5 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>64.5,-5.5,64.5,-1</points>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<intersection>-5.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>63,-5.5,63,-1</points>
<connection>
<GID>201</GID>
<name>OUT_0</name></connection>
<intersection>-5.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>76.5,-23,80,-23</points>
<connection>
<GID>208</GID>
<name>IN_0</name></connection>
<intersection>76.5 2</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>76.5,-9,79.5,-9</points>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<intersection>76.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-26,80,-26</points>
<intersection>55 3</intersection>
<intersection>63.5 6</intersection>
<intersection>65.5 5</intersection>
<intersection>80 7</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>55,-26,55,1.5</points>
<intersection>-26 1</intersection>
<intersection>1.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>55,1.5,79,1.5</points>
<connection>
<GID>204</GID>
<name>IN_1</name></connection>
<intersection>55 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>65.5,-26,65.5,-17.5</points>
<intersection>-26 1</intersection>
<intersection>-17.5 8</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>63.5,-26,63.5,-17.5</points>
<connection>
<GID>202</GID>
<name>OUT_0</name></connection>
<intersection>-26 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>80,-26,80,-25</points>
<connection>
<GID>208</GID>
<name>IN_1</name></connection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>65.5,-17.5,66,-17.5</points>
<connection>
<GID>197</GID>
<name>IN_0</name></connection>
<intersection>65.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-1,70.5,3.5</points>
<connection>
<GID>195</GID>
<name>OUT_0</name></connection>
<intersection>3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>70.5,3.5,79,3.5</points>
<connection>
<GID>204</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71.5,-17.5,71.5,-11</points>
<intersection>-17.5 2</intersection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71.5,-11,79.5,-11</points>
<connection>
<GID>206</GID>
<name>IN_1</name></connection>
<intersection>71.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71.5,-17.5,72,-17.5</points>
<connection>
<GID>197</GID>
<name>OUT_0</name></connection>
<intersection>71.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86,-24,87.5,-24</points>
<connection>
<GID>208</GID>
<name>OUT</name></connection>
<connection>
<GID>212</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,-10,87,-5.5</points>
<intersection>-10 2</intersection>
<intersection>-5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87,-5.5,88.5,-5.5</points>
<connection>
<GID>210</GID>
<name>IN_1</name></connection>
<intersection>87 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>85.5,-10,87,-10</points>
<connection>
<GID>206</GID>
<name>OUT</name></connection>
<intersection>87 0</intersection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86.5,-3.5,86.5,2.5</points>
<intersection>-3.5 1</intersection>
<intersection>2.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86.5,-3.5,88.5,-3.5</points>
<connection>
<GID>210</GID>
<name>IN_0</name></connection>
<intersection>86.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>85,2.5,86.5,2.5</points>
<connection>
<GID>204</GID>
<name>OUT</name></connection>
<intersection>86.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94.5,-4.5,95.5,-4.5</points>
<connection>
<GID>210</GID>
<name>OUT</name></connection>
<connection>
<GID>214</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33.5,-71.5,-33.5,-64.5</points>
<connection>
<GID>223</GID>
<name>IN_1</name></connection>
<connection>
<GID>223</GID>
<name>IN_0</name></connection>
<intersection>-70.5 1</intersection>
<intersection>-64.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-35.5,-70.5,-33.5,-70.5</points>
<connection>
<GID>233</GID>
<name>OUT_0</name></connection>
<intersection>-33.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-33.5,-64.5,-17.5,-64.5</points>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<intersection>-33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33.5,-87,-33.5,-79.5</points>
<connection>
<GID>224</GID>
<name>IN_1</name></connection>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<intersection>-86 1</intersection>
<intersection>-79.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-35,-86,-33.5,-86</points>
<connection>
<GID>234</GID>
<name>OUT_0</name></connection>
<intersection>-33.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-33.5,-79.5,-17,-79.5</points>
<connection>
<GID>226</GID>
<name>IN_1</name></connection>
<intersection>-33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-25,-93,-25,-66.5</points>
<intersection>-93 3</intersection>
<intersection>-86 2</intersection>
<intersection>-66.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-25,-66.5,-17.5,-66.5</points>
<connection>
<GID>225</GID>
<name>IN_1</name></connection>
<intersection>-25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-27.5,-86,-25,-86</points>
<connection>
<GID>224</GID>
<name>OUT</name></connection>
<intersection>-25 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-25,-93,-17,-93</points>
<connection>
<GID>227</GID>
<name>IN_1</name></connection>
<intersection>-25 0</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-27.5,-70.5,-20.5,-70.5</points>
<connection>
<GID>223</GID>
<name>OUT</name></connection>
<intersection>-20.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-20.5,-77.5,-20.5,-70.5</points>
<intersection>-77.5 4</intersection>
<intersection>-70.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-20.5,-77.5,-17,-77.5</points>
<connection>
<GID>226</GID>
<name>IN_0</name></connection>
<intersection>-20.5 3</intersection>
<intersection>-19.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-19.5,-91,-19.5,-77.5</points>
<intersection>-91 6</intersection>
<intersection>-77.5 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-19.5,-91,-17,-91</points>
<connection>
<GID>227</GID>
<name>IN_0</name></connection>
<intersection>-19.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5,-71,-5,-65.5</points>
<intersection>-71 1</intersection>
<intersection>-65.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-5,-71,1.5,-71</points>
<connection>
<GID>228</GID>
<name>IN_0</name></connection>
<intersection>-5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-11.5,-65.5,-5,-65.5</points>
<connection>
<GID>225</GID>
<name>OUT</name></connection>
<intersection>-5 0</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-78.5,-4.5,-73</points>
<intersection>-78.5 2</intersection>
<intersection>-73 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-73,1.5,-73</points>
<connection>
<GID>228</GID>
<name>IN_1</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-11,-78.5,-4.5,-78.5</points>
<connection>
<GID>226</GID>
<name>OUT</name></connection>
<intersection>-4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11,-92,-10,-92</points>
<connection>
<GID>236</GID>
<name>N_in0</name></connection>
<connection>
<GID>227</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7.5,-72,8.5,-72</points>
<connection>
<GID>238</GID>
<name>N_in0</name></connection>
<connection>
<GID>228</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 3>
<page 4>
<PageViewport>-71.6777,-209.554,218.783,-353.123</PageViewport>
<gate>
<ID>240</ID>
<type>AA_LABEL</type>
<position>42,9</position>
<gparam>LABEL_TEXT FULL ADDER USING AOI , NAND , NOR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>242</ID>
<type>AA_INVERTER</type>
<position>24.5,-22.5</position>
<input>
<ID>IN_0</ID>144 </input>
<output>
<ID>OUT_0</ID>148 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>243</ID>
<type>AA_INVERTER</type>
<position>24.5,-37</position>
<input>
<ID>IN_0</ID>145 </input>
<output>
<ID>OUT_0</ID>147 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>244</ID>
<type>AA_INVERTER</type>
<position>24.5,-52</position>
<input>
<ID>IN_0</ID>146 </input>
<output>
<ID>OUT_0</ID>159 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>246</ID>
<type>AA_LABEL</type>
<position>-7,-30</position>
<gparam>LABEL_TEXT AOI</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>248</ID>
<type>AA_TOGGLE</type>
<position>15,-22.5</position>
<output>
<ID>OUT_0</ID>144 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>249</ID>
<type>AA_TOGGLE</type>
<position>14.5,-37</position>
<output>
<ID>OUT_0</ID>145 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>250</ID>
<type>AA_TOGGLE</type>
<position>15.5,-52</position>
<output>
<ID>OUT_0</ID>146 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>252</ID>
<type>AA_AND3</type>
<position>61,-12</position>
<input>
<ID>IN_0</ID>144 </input>
<input>
<ID>IN_1</ID>147 </input>
<input>
<ID>IN_2</ID>146 </input>
<output>
<ID>OUT</ID>150 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>253</ID>
<type>AA_AND3</type>
<position>61,-21</position>
<input>
<ID>IN_0</ID>148 </input>
<input>
<ID>IN_1</ID>145 </input>
<input>
<ID>IN_2</ID>146 </input>
<output>
<ID>OUT</ID>151 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>254</ID>
<type>AA_AND3</type>
<position>61.5,-30</position>
<input>
<ID>IN_0</ID>144 </input>
<input>
<ID>IN_1</ID>145 </input>
<input>
<ID>IN_2</ID>159 </input>
<output>
<ID>OUT</ID>152 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>255</ID>
<type>AA_AND3</type>
<position>61.5,-39</position>
<input>
<ID>IN_0</ID>144 </input>
<input>
<ID>IN_1</ID>145 </input>
<input>
<ID>IN_2</ID>146 </input>
<output>
<ID>OUT</ID>153 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>256</ID>
<type>AA_AND3</type>
<position>61.5,-48</position>
<input>
<ID>IN_0</ID>148 </input>
<input>
<ID>IN_1</ID>147 </input>
<input>
<ID>IN_2</ID>146 </input>
<output>
<ID>OUT</ID>154 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>257</ID>
<type>AA_AND3</type>
<position>61.5,-57</position>
<input>
<ID>IN_0</ID>148 </input>
<input>
<ID>IN_1</ID>145 </input>
<input>
<ID>IN_2</ID>159 </input>
<output>
<ID>OUT</ID>155 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>258</ID>
<type>AA_AND3</type>
<position>61.5,-66</position>
<input>
<ID>IN_0</ID>144 </input>
<input>
<ID>IN_1</ID>147 </input>
<input>
<ID>IN_2</ID>159 </input>
<output>
<ID>OUT</ID>156 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>262</ID>
<type>AE_OR4</type>
<position>86,-24</position>
<input>
<ID>IN_0</ID>150 </input>
<input>
<ID>IN_1</ID>151 </input>
<input>
<ID>IN_2</ID>152 </input>
<input>
<ID>IN_3</ID>153 </input>
<output>
<ID>OUT</ID>157 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>263</ID>
<type>AE_OR4</type>
<position>86.5,-49</position>
<input>
<ID>IN_0</ID>153 </input>
<input>
<ID>IN_1</ID>154 </input>
<input>
<ID>IN_2</ID>155 </input>
<input>
<ID>IN_3</ID>156 </input>
<output>
<ID>OUT</ID>158 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>265</ID>
<type>AA_LABEL</type>
<position>129,-22.5</position>
<gparam>LABEL_TEXT CARRY : AB'C + A"BC + ABC' + ABC</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>266</ID>
<type>AA_LABEL</type>
<position>133,-47</position>
<gparam>LABEL_TEXT SUM : A'B'C + A'BC' + AB'C' + ABC</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>268</ID>
<type>GA_LED</type>
<position>92.5,-24</position>
<input>
<ID>N_in0</ID>157 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>269</ID>
<type>GA_LED</type>
<position>93,-49</position>
<input>
<ID>N_in0</ID>158 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>271</ID>
<type>AA_LABEL</type>
<position>-14,-145</position>
<gparam>LABEL_TEXT NAND</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>280</ID>
<type>BA_NAND2</type>
<position>5.5,-129.5</position>
<input>
<ID>IN_0</ID>161 </input>
<input>
<ID>IN_1</ID>161 </input>
<output>
<ID>OUT</ID>167 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>281</ID>
<type>BA_NAND2</type>
<position>6,-144.5</position>
<input>
<ID>IN_0</ID>162 </input>
<input>
<ID>IN_1</ID>162 </input>
<output>
<ID>OUT</ID>165 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>282</ID>
<type>BA_NAND2</type>
<position>6,-161</position>
<input>
<ID>IN_0</ID>163 </input>
<input>
<ID>IN_1</ID>163 </input>
<output>
<ID>OUT</ID>166 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>286</ID>
<type>AA_TOGGLE</type>
<position>-2,-129.5</position>
<output>
<ID>OUT_0</ID>161 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>287</ID>
<type>AA_TOGGLE</type>
<position>-2.5,-144.5</position>
<output>
<ID>OUT_0</ID>162 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>288</ID>
<type>AA_TOGGLE</type>
<position>-2,-161</position>
<output>
<ID>OUT_0</ID>163 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>292</ID>
<type>BA_NAND3</type>
<position>50,-112</position>
<input>
<ID>IN_0</ID>161 </input>
<input>
<ID>IN_1</ID>165 </input>
<input>
<ID>IN_2</ID>166 </input>
<output>
<ID>OUT</ID>169 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>293</ID>
<type>BA_NAND3</type>
<position>50,-123.5</position>
<input>
<ID>IN_0</ID>167 </input>
<input>
<ID>IN_1</ID>162 </input>
<input>
<ID>IN_2</ID>166 </input>
<output>
<ID>OUT</ID>170 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>294</ID>
<type>BA_NAND3</type>
<position>50,-134</position>
<input>
<ID>IN_0</ID>167 </input>
<input>
<ID>IN_1</ID>165 </input>
<input>
<ID>IN_2</ID>163 </input>
<output>
<ID>OUT</ID>171 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>295</ID>
<type>BA_NAND3</type>
<position>50.5,-144</position>
<input>
<ID>IN_0</ID>161 </input>
<input>
<ID>IN_1</ID>162 </input>
<input>
<ID>IN_2</ID>163 </input>
<output>
<ID>OUT</ID>172 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>296</ID>
<type>BA_NAND3</type>
<position>50.5,-154.5</position>
<input>
<ID>IN_0</ID>167 </input>
<input>
<ID>IN_1</ID>162 </input>
<input>
<ID>IN_2</ID>163 </input>
<output>
<ID>OUT</ID>173 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>297</ID>
<type>BA_NAND3</type>
<position>51,-166</position>
<input>
<ID>IN_0</ID>161 </input>
<input>
<ID>IN_1</ID>165 </input>
<input>
<ID>IN_2</ID>163 </input>
<output>
<ID>OUT</ID>174 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>298</ID>
<type>BA_NAND3</type>
<position>50.5,-176.5</position>
<input>
<ID>IN_0</ID>161 </input>
<input>
<ID>IN_1</ID>162 </input>
<input>
<ID>IN_2</ID>166 </input>
<output>
<ID>OUT</ID>175 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>301</ID>
<type>BA_NAND4</type>
<position>87.5,-123.5</position>
<input>
<ID>IN_0</ID>169 </input>
<input>
<ID>IN_1</ID>170 </input>
<input>
<ID>IN_2</ID>171 </input>
<input>
<ID>IN_3</ID>172 </input>
<output>
<ID>OUT</ID>176 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>302</ID>
<type>BA_NAND4</type>
<position>86.5,-154</position>
<input>
<ID>IN_0</ID>172 </input>
<input>
<ID>IN_1</ID>173 </input>
<input>
<ID>IN_2</ID>174 </input>
<input>
<ID>IN_3</ID>175 </input>
<output>
<ID>OUT</ID>177 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>303</ID>
<type>AA_LABEL</type>
<position>126.5,-124.5</position>
<gparam>LABEL_TEXT CARRY : AB'C + A"BC + ABC' + ABC</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>304</ID>
<type>AA_LABEL</type>
<position>125.5,-153.5</position>
<gparam>LABEL_TEXT SUM : A'B'C + A'BC' + AB'C' + ABC</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>306</ID>
<type>GA_LED</type>
<position>96.5,-123.5</position>
<input>
<ID>N_in0</ID>176 </input>
<input>
<ID>N_in3</ID>176 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>311</ID>
<type>GA_LED</type>
<position>94.5,-154.5</position>
<input>
<ID>N_in0</ID>177 </input>
<input>
<ID>N_in3</ID>177 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>312</ID>
<type>AA_LABEL</type>
<position>-22.5,-227.5</position>
<gparam>LABEL_TEXT NOR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>314</ID>
<type>BE_NOR3</type>
<position>60.5,-224</position>
<input>
<ID>IN_0</ID>178 </input>
<input>
<ID>IN_1</ID>179 </input>
<input>
<ID>IN_2</ID>183 </input>
<output>
<ID>OUT</ID>193 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>315</ID>
<type>BE_NOR3</type>
<position>61,-237.5</position>
<input>
<ID>IN_0</ID>184 </input>
<input>
<ID>IN_1</ID>179 </input>
<input>
<ID>IN_2</ID>180 </input>
<output>
<ID>OUT</ID>194 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>316</ID>
<type>BE_NOR3</type>
<position>61,-251.5</position>
<input>
<ID>IN_0</ID>178 </input>
<input>
<ID>IN_1</ID>185 </input>
<input>
<ID>IN_2</ID>180 </input>
<output>
<ID>OUT</ID>195 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>317</ID>
<type>BE_NOR3</type>
<position>61.5,-265</position>
<input>
<ID>IN_0</ID>184 </input>
<input>
<ID>IN_1</ID>185 </input>
<input>
<ID>IN_2</ID>183 </input>
<output>
<ID>OUT</ID>196 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>318</ID>
<type>BE_NOR3</type>
<position>62,-277.5</position>
<input>
<ID>IN_0</ID>178 </input>
<input>
<ID>IN_1</ID>185 </input>
<input>
<ID>IN_2</ID>183 </input>
<output>
<ID>OUT</ID>197 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>319</ID>
<type>BE_NOR3</type>
<position>62.5,-290</position>
<input>
<ID>IN_0</ID>184 </input>
<input>
<ID>IN_1</ID>180 </input>
<input>
<ID>IN_2</ID>183 </input>
<output>
<ID>OUT</ID>198 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>320</ID>
<type>BE_NOR3</type>
<position>62.5,-303.5</position>
<input>
<ID>IN_0</ID>184 </input>
<input>
<ID>IN_1</ID>185 </input>
<input>
<ID>IN_2</ID>180 </input>
<output>
<ID>OUT</ID>199 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>326</ID>
<type>BE_NOR2</type>
<position>21,-235.5</position>
<input>
<ID>IN_0</ID>178 </input>
<input>
<ID>IN_1</ID>178 </input>
<output>
<ID>OUT</ID>184 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>327</ID>
<type>BE_NOR2</type>
<position>21,-259.5</position>
<input>
<ID>IN_0</ID>179 </input>
<input>
<ID>IN_1</ID>179 </input>
<output>
<ID>OUT</ID>185 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>328</ID>
<type>BE_NOR2</type>
<position>22,-284.5</position>
<input>
<ID>IN_0</ID>180 </input>
<input>
<ID>IN_1</ID>180 </input>
<output>
<ID>OUT</ID>183 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>330</ID>
<type>AA_TOGGLE</type>
<position>8.5,-235.5</position>
<output>
<ID>OUT_0</ID>178 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>331</ID>
<type>AA_TOGGLE</type>
<position>9,-259.5</position>
<output>
<ID>OUT_0</ID>179 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>332</ID>
<type>AA_TOGGLE</type>
<position>9.5,-285</position>
<output>
<ID>OUT_0</ID>180 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>336</ID>
<type>GA_LED</type>
<position>107.5,-240.5</position>
<input>
<ID>N_in0</ID>201 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>338</ID>
<type>GA_LED</type>
<position>110.5,-291</position>
<input>
<ID>N_in0</ID>200 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>339</ID>
<type>AA_LABEL</type>
<position>138,-240.5</position>
<gparam>LABEL_TEXT CARRY : AB'C + A"BC + ABC' + ABC</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>340</ID>
<type>AA_LABEL</type>
<position>139,-290.5</position>
<gparam>LABEL_TEXT SUM : A'B'C + A'BC' + AB'C' + ABC</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>344</ID>
<type>BE_NOR4</type>
<position>93.5,-233</position>
<input>
<ID>IN_0</ID>193 </input>
<input>
<ID>IN_1</ID>194 </input>
<input>
<ID>IN_2</ID>195 </input>
<input>
<ID>IN_3</ID>196 </input>
<output>
<ID>OUT</ID>201 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>345</ID>
<type>BE_NOR4</type>
<position>95,-291.5</position>
<input>
<ID>IN_0</ID>196 </input>
<input>
<ID>IN_1</ID>197 </input>
<input>
<ID>IN_2</ID>198 </input>
<input>
<ID>IN_3</ID>199 </input>
<output>
<ID>OUT</ID>200 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<wire>
<ID>193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77,-230,77,-224</points>
<intersection>-230 1</intersection>
<intersection>-224 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77,-230,90.5,-230</points>
<connection>
<GID>344</GID>
<name>IN_0</name></connection>
<intersection>77 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-224,77,-224</points>
<connection>
<GID>314</GID>
<name>OUT</name></connection>
<intersection>77 0</intersection></hsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77,-237.5,77,-232</points>
<intersection>-237.5 2</intersection>
<intersection>-232 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77,-232,90.5,-232</points>
<connection>
<GID>344</GID>
<name>IN_1</name></connection>
<intersection>77 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>64,-237.5,77,-237.5</points>
<connection>
<GID>315</GID>
<name>OUT</name></connection>
<intersection>77 0</intersection></hsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-251.5,74.5,-230.5</points>
<intersection>-251.5 2</intersection>
<intersection>-230.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,-230.5,90.5,-230.5</points>
<intersection>74.5 0</intersection>
<intersection>90.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>64,-251.5,74.5,-251.5</points>
<connection>
<GID>316</GID>
<name>OUT</name></connection>
<intersection>74.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>90.5,-234,90.5,-230.5</points>
<connection>
<GID>344</GID>
<name>IN_2</name></connection>
<intersection>-230.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-288.5,77.5,-236</points>
<intersection>-288.5 3</intersection>
<intersection>-265 2</intersection>
<intersection>-236 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77.5,-236,90.5,-236</points>
<connection>
<GID>344</GID>
<name>IN_3</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>64.5,-265,77.5,-265</points>
<connection>
<GID>317</GID>
<name>OUT</name></connection>
<intersection>77.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>77.5,-288.5,92,-288.5</points>
<connection>
<GID>345</GID>
<name>IN_0</name></connection>
<intersection>77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78.5,-290.5,78.5,-277.5</points>
<intersection>-290.5 2</intersection>
<intersection>-277.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65,-277.5,78.5,-277.5</points>
<connection>
<GID>318</GID>
<name>OUT</name></connection>
<intersection>78.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>78.5,-290.5,92,-290.5</points>
<connection>
<GID>345</GID>
<name>IN_1</name></connection>
<intersection>78.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>65.5,-292.5,92,-292.5</points>
<connection>
<GID>345</GID>
<name>IN_2</name></connection>
<intersection>65.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>65.5,-292.5,65.5,-290</points>
<connection>
<GID>319</GID>
<name>OUT</name></connection>
<intersection>-292.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78.5,-303.5,78.5,-294.5</points>
<intersection>-303.5 1</intersection>
<intersection>-294.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65.5,-303.5,78.5,-303.5</points>
<connection>
<GID>320</GID>
<name>OUT</name></connection>
<intersection>78.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>78.5,-294.5,92,-294.5</points>
<connection>
<GID>345</GID>
<name>IN_3</name></connection>
<intersection>78.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,-291.5,104,-291</points>
<intersection>-291.5 2</intersection>
<intersection>-291 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104,-291,109.5,-291</points>
<connection>
<GID>338</GID>
<name>N_in0</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>99,-291.5,104,-291.5</points>
<connection>
<GID>345</GID>
<name>OUT</name></connection>
<intersection>104 0</intersection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,-240.5,102,-233</points>
<intersection>-240.5 1</intersection>
<intersection>-233 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>102,-240.5,106.5,-240.5</points>
<connection>
<GID>336</GID>
<name>N_in0</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-233,102,-233</points>
<connection>
<GID>344</GID>
<name>OUT</name></connection>
<intersection>102 0</intersection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17,-22.5,21.5,-22.5</points>
<connection>
<GID>248</GID>
<name>OUT_0</name></connection>
<connection>
<GID>242</GID>
<name>IN_0</name></connection>
<intersection>20 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>20,-22.5,20,-10</points>
<intersection>-22.5 1</intersection>
<intersection>-10 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>20,-10,58,-10</points>
<connection>
<GID>252</GID>
<name>IN_0</name></connection>
<intersection>20 3</intersection>
<intersection>52.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>52.5,-28,52.5,-10</points>
<intersection>-28 6</intersection>
<intersection>-10 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>52.5,-28,58.5,-28</points>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<intersection>52.5 5</intersection>
<intersection>56 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>56,-37,56,-28</points>
<intersection>-37 9</intersection>
<intersection>-28 6</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>40.5,-37,58.5,-37</points>
<connection>
<GID>255</GID>
<name>IN_0</name></connection>
<intersection>40.5 11</intersection>
<intersection>56 8</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>40.5,-64,40.5,-37</points>
<intersection>-64 12</intersection>
<intersection>-37 9</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>40.5,-64,58.5,-64</points>
<connection>
<GID>258</GID>
<name>IN_0</name></connection>
<intersection>40.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-37,21.5,-37</points>
<connection>
<GID>243</GID>
<name>IN_0</name></connection>
<connection>
<GID>249</GID>
<name>OUT_0</name></connection>
<intersection>20.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>20.5,-37,20.5,-20</points>
<intersection>-37 1</intersection>
<intersection>-20 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>20.5,-20,50.5,-20</points>
<intersection>20.5 3</intersection>
<intersection>50.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>50.5,-30,50.5,-20</points>
<intersection>-30 6</intersection>
<intersection>-21 7</intersection>
<intersection>-20 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>50.5,-30,58.5,-30</points>
<connection>
<GID>254</GID>
<name>IN_1</name></connection>
<intersection>50.5 5</intersection>
<intersection>58 8</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>50.5,-21,58,-21</points>
<connection>
<GID>253</GID>
<name>IN_1</name></connection>
<intersection>50.5 5</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>58,-39,58,-30</points>
<intersection>-39 9</intersection>
<intersection>-30 6</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>38.5,-39,58.5,-39</points>
<connection>
<GID>255</GID>
<name>IN_1</name></connection>
<intersection>38.5 10</intersection>
<intersection>58 8</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>38.5,-57,38.5,-39</points>
<intersection>-57 11</intersection>
<intersection>-39 9</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>38.5,-57,58.5,-57</points>
<connection>
<GID>257</GID>
<name>IN_1</name></connection>
<intersection>38.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17.5,-56,29.5,-56</points>
<intersection>17.5 8</intersection>
<intersection>21.5 7</intersection>
<intersection>29.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>29.5,-56,29.5,-14</points>
<intersection>-56 1</intersection>
<intersection>-25 6</intersection>
<intersection>-14 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>29.5,-14,58,-14</points>
<connection>
<GID>252</GID>
<name>IN_2</name></connection>
<intersection>29.5 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>29.5,-25,58,-25</points>
<intersection>29.5 4</intersection>
<intersection>46.5 10</intersection>
<intersection>58 9</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>21.5,-56,21.5,-52</points>
<connection>
<GID>244</GID>
<name>IN_0</name></connection>
<intersection>-56 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>17.5,-56,17.5,-52</points>
<intersection>-56 1</intersection>
<intersection>-52 13</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>58,-25,58,-23</points>
<connection>
<GID>253</GID>
<name>IN_2</name></connection>
<intersection>-25 6</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>46.5,-41,46.5,-25</points>
<intersection>-41 11</intersection>
<intersection>-25 6</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>46.5,-41,58.5,-41</points>
<connection>
<GID>255</GID>
<name>IN_2</name></connection>
<intersection>46.5 10</intersection>
<intersection>58.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>58.5,-50,58.5,-41</points>
<connection>
<GID>256</GID>
<name>IN_2</name></connection>
<intersection>-41 11</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>17.5,-52,17.5,-52</points>
<connection>
<GID>250</GID>
<name>OUT_0</name></connection>
<intersection>17.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-48,32.5,-12</points>
<intersection>-48 3</intersection>
<intersection>-37 1</intersection>
<intersection>-12 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-37,32.5,-37</points>
<connection>
<GID>243</GID>
<name>OUT_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-12,58,-12</points>
<connection>
<GID>252</GID>
<name>IN_1</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>32.5,-48,58.5,-48</points>
<connection>
<GID>256</GID>
<name>IN_1</name></connection>
<intersection>32.5 0</intersection>
<intersection>43.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>43.5,-66,43.5,-48</points>
<intersection>-66 5</intersection>
<intersection>-48 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>43.5,-66,58.5,-66</points>
<connection>
<GID>258</GID>
<name>IN_1</name></connection>
<intersection>43.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-22.5,32.5,-19</points>
<intersection>-22.5 3</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-19,58,-19</points>
<connection>
<GID>253</GID>
<name>IN_0</name></connection>
<intersection>32.5 0</intersection>
<intersection>43.5 4</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>27.5,-22.5,32.5,-22.5</points>
<connection>
<GID>242</GID>
<name>OUT_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>43.5,-46,43.5,-19</points>
<intersection>-46 5</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>43.5,-46,58.5,-46</points>
<connection>
<GID>256</GID>
<name>IN_0</name></connection>
<intersection>43.5 4</intersection>
<intersection>56 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>56,-55,56,-46</points>
<intersection>-55 7</intersection>
<intersection>-46 5</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>56,-55,58.5,-55</points>
<connection>
<GID>257</GID>
<name>IN_0</name></connection>
<intersection>56 6</intersection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-18.5,73.5,-12</points>
<intersection>-18.5 1</intersection>
<intersection>-12 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73.5,-18.5,83,-18.5</points>
<intersection>73.5 0</intersection>
<intersection>83 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>64,-12,73.5,-12</points>
<connection>
<GID>252</GID>
<name>OUT</name></connection>
<intersection>73.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>83,-21,83,-18.5</points>
<connection>
<GID>262</GID>
<name>IN_0</name></connection>
<intersection>-18.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-23,73.5,-21</points>
<intersection>-23 1</intersection>
<intersection>-21 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73.5,-23,83,-23</points>
<connection>
<GID>262</GID>
<name>IN_1</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>64,-21,73.5,-21</points>
<connection>
<GID>253</GID>
<name>OUT</name></connection>
<intersection>73.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-30,73.5,-25</points>
<intersection>-30 2</intersection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73.5,-25,83,-25</points>
<connection>
<GID>262</GID>
<name>IN_2</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>64.5,-30,73.5,-30</points>
<connection>
<GID>254</GID>
<name>OUT</name></connection>
<intersection>73.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-46,76.5,-27</points>
<intersection>-46 3</intersection>
<intersection>-39 2</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76.5,-27,83,-27</points>
<connection>
<GID>262</GID>
<name>IN_3</name></connection>
<intersection>76.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>64.5,-39,76.5,-39</points>
<connection>
<GID>255</GID>
<name>OUT</name></connection>
<intersection>76.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>76.5,-46,83.5,-46</points>
<connection>
<GID>263</GID>
<name>IN_0</name></connection>
<intersection>76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64.5,-48,83.5,-48</points>
<connection>
<GID>256</GID>
<name>OUT</name></connection>
<connection>
<GID>263</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,-57,74,-50</points>
<intersection>-57 1</intersection>
<intersection>-50 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64.5,-57,74,-57</points>
<connection>
<GID>257</GID>
<name>OUT</name></connection>
<intersection>74 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>74,-50,83.5,-50</points>
<connection>
<GID>263</GID>
<name>IN_2</name></connection>
<intersection>74 0</intersection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-66,76.5,-52</points>
<intersection>-66 1</intersection>
<intersection>-52 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64.5,-66,76.5,-66</points>
<connection>
<GID>258</GID>
<name>OUT</name></connection>
<intersection>76.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>76.5,-52,83.5,-52</points>
<connection>
<GID>263</GID>
<name>IN_3</name></connection>
<intersection>76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90,-24,91.5,-24</points>
<connection>
<GID>268</GID>
<name>N_in0</name></connection>
<connection>
<GID>262</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90.5,-49,92,-49</points>
<connection>
<GID>269</GID>
<name>N_in0</name></connection>
<intersection>90.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>90.5,-49,90.5,-49</points>
<connection>
<GID>263</GID>
<name>OUT</name></connection>
<intersection>-49 1</intersection></vsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,-59,41.5,-32</points>
<intersection>-59 2</intersection>
<intersection>-52 1</intersection>
<intersection>-32 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-52,41.5,-52</points>
<connection>
<GID>244</GID>
<name>OUT_0</name></connection>
<intersection>41.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>41.5,-59,58.5,-59</points>
<connection>
<GID>257</GID>
<name>IN_2</name></connection>
<intersection>41.5 0</intersection>
<intersection>58.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>58.5,-68,58.5,-59</points>
<connection>
<GID>258</GID>
<name>IN_2</name></connection>
<intersection>-59 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>41.5,-32,58.5,-32</points>
<connection>
<GID>254</GID>
<name>IN_2</name></connection>
<intersection>41.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.5,-130.5,2.5,-110</points>
<connection>
<GID>280</GID>
<name>IN_1</name></connection>
<connection>
<GID>280</GID>
<name>IN_0</name></connection>
<intersection>-129.5 1</intersection>
<intersection>-110 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0,-129.5,2.5,-129.5</points>
<connection>
<GID>286</GID>
<name>OUT_0</name></connection>
<intersection>2.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>2.5,-110,47,-110</points>
<connection>
<GID>292</GID>
<name>IN_0</name></connection>
<intersection>2.5 0</intersection>
<intersection>40.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>40.5,-142,40.5,-110</points>
<intersection>-142 7</intersection>
<intersection>-110 3</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>27.5,-142,47.5,-142</points>
<connection>
<GID>295</GID>
<name>IN_0</name></connection>
<intersection>27.5 8</intersection>
<intersection>40.5 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>27.5,-174.5,27.5,-142</points>
<intersection>-174.5 9</intersection>
<intersection>-164 10</intersection>
<intersection>-142 7</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>27.5,-174.5,47.5,-174.5</points>
<connection>
<GID>298</GID>
<name>IN_0</name></connection>
<intersection>27.5 8</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>27.5,-164,48,-164</points>
<connection>
<GID>297</GID>
<name>IN_0</name></connection>
<intersection>27.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-145.5,3,-123.5</points>
<connection>
<GID>281</GID>
<name>IN_1</name></connection>
<connection>
<GID>281</GID>
<name>IN_0</name></connection>
<intersection>-144.5 1</intersection>
<intersection>-123.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-0.5,-144.5,3,-144.5</points>
<connection>
<GID>287</GID>
<name>OUT_0</name></connection>
<intersection>3 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>3,-123.5,47,-123.5</points>
<connection>
<GID>293</GID>
<name>IN_1</name></connection>
<intersection>3 0</intersection>
<intersection>44 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>44,-144.5,44,-123.5</points>
<intersection>-144.5 4</intersection>
<intersection>-123.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>42.5,-144.5,47.5,-144.5</points>
<intersection>42.5 6</intersection>
<intersection>44 3</intersection>
<intersection>47.5 8</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>42.5,-154.5,42.5,-144.5</points>
<intersection>-154.5 7</intersection>
<intersection>-144.5 4</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>38.5,-154.5,47.5,-154.5</points>
<connection>
<GID>296</GID>
<name>IN_1</name></connection>
<intersection>38.5 9</intersection>
<intersection>42.5 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>47.5,-144.5,47.5,-144</points>
<connection>
<GID>295</GID>
<name>IN_1</name></connection>
<intersection>-144.5 4</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>38.5,-176.5,38.5,-154.5</points>
<intersection>-176.5 10</intersection>
<intersection>-154.5 7</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>38.5,-176.5,47.5,-176.5</points>
<connection>
<GID>298</GID>
<name>IN_1</name></connection>
<intersection>38.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1.5,-162,1.5,-136</points>
<intersection>-162 3</intersection>
<intersection>-161 1</intersection>
<intersection>-160 4</intersection>
<intersection>-136 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0,-161,1.5,-161</points>
<connection>
<GID>288</GID>
<name>OUT_0</name></connection>
<intersection>1.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1.5,-136,47,-136</points>
<connection>
<GID>294</GID>
<name>IN_2</name></connection>
<intersection>1.5 0</intersection>
<intersection>33 5</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>1.5,-162,3,-162</points>
<connection>
<GID>282</GID>
<name>IN_1</name></connection>
<intersection>1.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>1.5,-160,3,-160</points>
<connection>
<GID>282</GID>
<name>IN_0</name></connection>
<intersection>1.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>33,-146,33,-136</points>
<intersection>-146 6</intersection>
<intersection>-136 2</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>33,-146,47.5,-146</points>
<connection>
<GID>295</GID>
<name>IN_2</name></connection>
<intersection>33 5</intersection>
<intersection>41 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>41,-156.5,41,-146</points>
<intersection>-156.5 8</intersection>
<intersection>-146 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>33,-156.5,47.5,-156.5</points>
<connection>
<GID>296</GID>
<name>IN_2</name></connection>
<intersection>33 9</intersection>
<intersection>41 7</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>33,-168,33,-156.5</points>
<intersection>-168 10</intersection>
<intersection>-156.5 8</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>33,-168,48,-168</points>
<connection>
<GID>297</GID>
<name>IN_2</name></connection>
<intersection>33 9</intersection></hsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-144.5,23.5,-112</points>
<intersection>-144.5 1</intersection>
<intersection>-134 3</intersection>
<intersection>-112 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-144.5,23.5,-144.5</points>
<connection>
<GID>281</GID>
<name>OUT</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23.5,-112,47,-112</points>
<connection>
<GID>292</GID>
<name>IN_1</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>23.5,-134,47,-134</points>
<connection>
<GID>294</GID>
<name>IN_1</name></connection>
<intersection>23.5 0</intersection>
<intersection>45 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>45,-166,45,-134</points>
<intersection>-166 5</intersection>
<intersection>-134 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>45,-166,48,-166</points>
<connection>
<GID>297</GID>
<name>IN_1</name></connection>
<intersection>45 4</intersection></hsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,-178.5,18.5,-114</points>
<intersection>-178.5 6</intersection>
<intersection>-161 1</intersection>
<intersection>-114 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-161,18.5,-161</points>
<connection>
<GID>282</GID>
<name>OUT</name></connection>
<intersection>18.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18.5,-114,47,-114</points>
<connection>
<GID>292</GID>
<name>IN_2</name></connection>
<intersection>18.5 0</intersection>
<intersection>45 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>45,-125.5,45,-114</points>
<intersection>-125.5 4</intersection>
<intersection>-114 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>45,-125.5,47,-125.5</points>
<connection>
<GID>293</GID>
<name>IN_2</name></connection>
<intersection>45 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>18.5,-178.5,47.5,-178.5</points>
<connection>
<GID>298</GID>
<name>IN_2</name></connection>
<intersection>18.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-129.5,27.5,-121.5</points>
<intersection>-129.5 2</intersection>
<intersection>-121.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-121.5,47,-121.5</points>
<connection>
<GID>293</GID>
<name>IN_0</name></connection>
<intersection>27.5 0</intersection>
<intersection>47 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-129.5,27.5,-129.5</points>
<connection>
<GID>280</GID>
<name>OUT</name></connection>
<intersection>27.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>47,-152.5,47,-121.5</points>
<connection>
<GID>294</GID>
<name>IN_0</name></connection>
<intersection>-152.5 5</intersection>
<intersection>-121.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>47,-152.5,47.5,-152.5</points>
<connection>
<GID>296</GID>
<name>IN_0</name></connection>
<intersection>47 3</intersection></hsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-120.5,68.5,-112</points>
<intersection>-120.5 1</intersection>
<intersection>-112 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-120.5,84.5,-120.5</points>
<connection>
<GID>301</GID>
<name>IN_0</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53,-112,68.5,-112</points>
<connection>
<GID>292</GID>
<name>OUT</name></connection>
<intersection>68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-122.5,84.5,-122.5</points>
<connection>
<GID>301</GID>
<name>IN_1</name></connection>
<intersection>53 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>53,-123.5,53,-122.5</points>
<connection>
<GID>293</GID>
<name>OUT</name></connection>
<intersection>-122.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-134,68.5,-124.5</points>
<intersection>-134 2</intersection>
<intersection>-124.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-124.5,84.5,-124.5</points>
<connection>
<GID>301</GID>
<name>IN_2</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53,-134,68.5,-134</points>
<connection>
<GID>294</GID>
<name>OUT</name></connection>
<intersection>68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71,-151,71,-126.5</points>
<intersection>-151 3</intersection>
<intersection>-144 2</intersection>
<intersection>-126.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71,-126.5,84.5,-126.5</points>
<connection>
<GID>301</GID>
<name>IN_3</name></connection>
<intersection>71 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53.5,-144,71,-144</points>
<connection>
<GID>295</GID>
<name>OUT</name></connection>
<intersection>71 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>71,-151,83.5,-151</points>
<connection>
<GID>302</GID>
<name>IN_0</name></connection>
<intersection>71 0</intersection></hsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53.5,-153,83.5,-153</points>
<connection>
<GID>302</GID>
<name>IN_1</name></connection>
<intersection>53.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>53.5,-154.5,53.5,-153</points>
<connection>
<GID>296</GID>
<name>OUT</name></connection>
<intersection>-153 1</intersection></vsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-166,68.5,-155</points>
<intersection>-166 2</intersection>
<intersection>-155 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-155,83.5,-155</points>
<connection>
<GID>302</GID>
<name>IN_2</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54,-166,68.5,-166</points>
<connection>
<GID>297</GID>
<name>OUT</name></connection>
<intersection>68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,-176.5,72.5,-157</points>
<intersection>-176.5 2</intersection>
<intersection>-157 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72.5,-157,83.5,-157</points>
<connection>
<GID>302</GID>
<name>IN_3</name></connection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53.5,-176.5,72.5,-176.5</points>
<connection>
<GID>298</GID>
<name>OUT</name></connection>
<intersection>72.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90.5,-123.5,96.5,-123.5</points>
<connection>
<GID>301</GID>
<name>OUT</name></connection>
<connection>
<GID>306</GID>
<name>N_in0</name></connection>
<intersection>96.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>96.5,-123.5,96.5,-122.5</points>
<connection>
<GID>306</GID>
<name>N_in3</name></connection>
<intersection>-123.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>89.5,-154.5,94.5,-154.5</points>
<connection>
<GID>311</GID>
<name>N_in0</name></connection>
<intersection>89.5 4</intersection>
<intersection>94.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>94.5,-154.5,94.5,-153.5</points>
<connection>
<GID>311</GID>
<name>N_in3</name></connection>
<intersection>-154.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>89.5,-154.5,89.5,-154</points>
<connection>
<GID>302</GID>
<name>OUT</name></connection>
<intersection>-154.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-236.5,18,-222</points>
<connection>
<GID>326</GID>
<name>IN_1</name></connection>
<connection>
<GID>326</GID>
<name>IN_0</name></connection>
<intersection>-235.5 1</intersection>
<intersection>-222 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10.5,-235.5,18,-235.5</points>
<connection>
<GID>330</GID>
<name>OUT_0</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18,-222,58,-222</points>
<connection>
<GID>314</GID>
<name>IN_0</name></connection>
<intersection>18 0</intersection>
<intersection>58 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>58,-275.5,58,-222</points>
<connection>
<GID>316</GID>
<name>IN_0</name></connection>
<intersection>-275.5 5</intersection>
<intersection>-222 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>58,-275.5,59,-275.5</points>
<connection>
<GID>318</GID>
<name>IN_0</name></connection>
<intersection>58 3</intersection></hsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15.5,-260.5,15.5,-224</points>
<intersection>-260.5 3</intersection>
<intersection>-259.5 1</intersection>
<intersection>-258.5 4</intersection>
<intersection>-224 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11,-259.5,15.5,-259.5</points>
<connection>
<GID>331</GID>
<name>OUT_0</name></connection>
<intersection>15.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15.5,-224,57.5,-224</points>
<connection>
<GID>314</GID>
<name>IN_1</name></connection>
<intersection>15.5 0</intersection>
<intersection>53.5 5</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>15.5,-260.5,18,-260.5</points>
<connection>
<GID>327</GID>
<name>IN_1</name></connection>
<intersection>15.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>15.5,-258.5,18,-258.5</points>
<connection>
<GID>327</GID>
<name>IN_0</name></connection>
<intersection>15.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>53.5,-237.5,53.5,-224</points>
<intersection>-237.5 6</intersection>
<intersection>-224 2</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>53.5,-237.5,58,-237.5</points>
<connection>
<GID>315</GID>
<name>IN_1</name></connection>
<intersection>53.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-285.5,17.5,-239.5</points>
<intersection>-285.5 3</intersection>
<intersection>-285 1</intersection>
<intersection>-283.5 4</intersection>
<intersection>-239.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11.5,-285,17.5,-285</points>
<connection>
<GID>332</GID>
<name>OUT_0</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17.5,-239.5,58,-239.5</points>
<connection>
<GID>315</GID>
<name>IN_2</name></connection>
<intersection>17.5 0</intersection>
<intersection>50.5 5</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>17.5,-285.5,19,-285.5</points>
<connection>
<GID>328</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>17.5,-283.5,19,-283.5</points>
<connection>
<GID>328</GID>
<name>IN_0</name></connection>
<intersection>17.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>50.5,-253.5,50.5,-239.5</points>
<intersection>-253.5 6</intersection>
<intersection>-239.5 2</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>50.5,-253.5,58,-253.5</points>
<connection>
<GID>316</GID>
<name>IN_2</name></connection>
<intersection>50.5 5</intersection>
<intersection>56 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>56,-290,56,-253.5</points>
<intersection>-290 8</intersection>
<intersection>-253.5 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>55,-290,59.5,-290</points>
<connection>
<GID>319</GID>
<name>IN_1</name></connection>
<intersection>55 9</intersection>
<intersection>56 7</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>55,-305.5,55,-290</points>
<intersection>-305.5 10</intersection>
<intersection>-290 8</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>55,-305.5,59.5,-305.5</points>
<connection>
<GID>320</GID>
<name>IN_2</name></connection>
<intersection>55 9</intersection></hsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-284.5,38,-226</points>
<intersection>-284.5 1</intersection>
<intersection>-267 4</intersection>
<intersection>-226 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-284.5,38,-284.5</points>
<connection>
<GID>328</GID>
<name>OUT</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38,-226,57.5,-226</points>
<connection>
<GID>314</GID>
<name>IN_2</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>38,-267,58.5,-267</points>
<connection>
<GID>317</GID>
<name>IN_2</name></connection>
<intersection>38 0</intersection>
<intersection>49.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>49.5,-279.5,49.5,-267</points>
<intersection>-279.5 6</intersection>
<intersection>-267 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>49.5,-279.5,59,-279.5</points>
<connection>
<GID>318</GID>
<name>IN_2</name></connection>
<intersection>49.5 5</intersection>
<intersection>54 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>54,-292,54,-279.5</points>
<intersection>-292 8</intersection>
<intersection>-279.5 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>54,-292,59.5,-292</points>
<connection>
<GID>319</GID>
<name>IN_2</name></connection>
<intersection>54 7</intersection></hsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24,-235.5,58,-235.5</points>
<connection>
<GID>326</GID>
<name>OUT</name></connection>
<connection>
<GID>315</GID>
<name>IN_0</name></connection>
<intersection>57 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>57,-288,57,-235.5</points>
<intersection>-288 4</intersection>
<intersection>-263 5</intersection>
<intersection>-235.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>57,-288,59.5,-288</points>
<connection>
<GID>319</GID>
<name>IN_0</name></connection>
<intersection>57 3</intersection>
<intersection>59.5 6</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>57,-263,58.5,-263</points>
<connection>
<GID>317</GID>
<name>IN_0</name></connection>
<intersection>57 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>59.5,-301.5,59.5,-288</points>
<connection>
<GID>320</GID>
<name>IN_0</name></connection>
<intersection>-288 4</intersection></vsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,-259.5,41,-251.5</points>
<intersection>-259.5 1</intersection>
<intersection>-251.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24,-259.5,41,-259.5</points>
<connection>
<GID>327</GID>
<name>OUT</name></connection>
<intersection>41 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>41,-251.5,58,-251.5</points>
<connection>
<GID>316</GID>
<name>IN_1</name></connection>
<intersection>41 0</intersection>
<intersection>45.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>45.5,-265,45.5,-251.5</points>
<intersection>-265 4</intersection>
<intersection>-251.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>45.5,-265,58.5,-265</points>
<connection>
<GID>317</GID>
<name>IN_1</name></connection>
<intersection>45.5 3</intersection>
<intersection>53 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>53,-277.5,53,-265</points>
<intersection>-277.5 6</intersection>
<intersection>-265 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>46,-277.5,59,-277.5</points>
<connection>
<GID>318</GID>
<name>IN_1</name></connection>
<intersection>46 7</intersection>
<intersection>53 5</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>46,-303.5,46,-277.5</points>
<intersection>-303.5 8</intersection>
<intersection>-277.5 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>46,-303.5,59.5,-303.5</points>
<connection>
<GID>320</GID>
<name>IN_1</name></connection>
<intersection>46 7</intersection></hsegment></shape></wire></page 4>
<page 5>
<PageViewport>-20.4,-38.8222,142.8,-119.489</PageViewport>
<gate>
<ID>342</ID>
<type>AA_LABEL</type>
<position>32.5,16.5</position>
<gparam>LABEL_TEXT SUBTRACTOR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>347</ID>
<type>AA_INVERTER</type>
<position>22,-8</position>
<input>
<ID>IN_0</ID>204 </input>
<output>
<ID>OUT_0</ID>202 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>348</ID>
<type>AA_INVERTER</type>
<position>22,-27</position>
<input>
<ID>IN_0</ID>203 </input>
<output>
<ID>OUT_0</ID>205 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>351</ID>
<type>AA_AND2</type>
<position>43,-2</position>
<input>
<ID>IN_0</ID>202 </input>
<input>
<ID>IN_1</ID>203 </input>
<output>
<ID>OUT</ID>206 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>352</ID>
<type>AA_AND2</type>
<position>43.5,-17.5</position>
<input>
<ID>IN_0</ID>204 </input>
<input>
<ID>IN_1</ID>205 </input>
<output>
<ID>OUT</ID>207 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>353</ID>
<type>AA_AND2</type>
<position>43,-36</position>
<input>
<ID>IN_0</ID>202 </input>
<input>
<ID>IN_1</ID>203 </input>
<output>
<ID>OUT</ID>209 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>355</ID>
<type>AE_OR2</type>
<position>58,-9.5</position>
<input>
<ID>IN_0</ID>206 </input>
<input>
<ID>IN_1</ID>207 </input>
<output>
<ID>OUT</ID>208 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>357</ID>
<type>AA_TOGGLE</type>
<position>3.5,-9.5</position>
<output>
<ID>OUT_0</ID>204 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>358</ID>
<type>AA_TOGGLE</type>
<position>4.5,-27</position>
<output>
<ID>OUT_0</ID>203 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>360</ID>
<type>GA_LED</type>
<position>64.5,-9.5</position>
<input>
<ID>N_in0</ID>208 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>361</ID>
<type>GA_LED</type>
<position>49,-36.5</position>
<input>
<ID>N_in0</ID>209 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>364</ID>
<type>AA_TOGGLE</type>
<position>-3,-75.5</position>
<output>
<ID>OUT_0</ID>222 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>365</ID>
<type>AA_TOGGLE</type>
<position>-1,-94</position>
<output>
<ID>OUT_0</ID>215 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>371</ID>
<type>BA_NAND2</type>
<position>18.5,-75.5</position>
<input>
<ID>IN_0</ID>222 </input>
<input>
<ID>IN_1</ID>222 </input>
<output>
<ID>OUT</ID>216 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>372</ID>
<type>BA_NAND2</type>
<position>17,-93.5</position>
<input>
<ID>IN_0</ID>215 </input>
<input>
<ID>IN_1</ID>215 </input>
<output>
<ID>OUT</ID>217 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>374</ID>
<type>BA_NAND2</type>
<position>41.5,-74.5</position>
<input>
<ID>IN_0</ID>216 </input>
<input>
<ID>IN_1</ID>215 </input>
<output>
<ID>OUT</ID>218 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>375</ID>
<type>BA_NAND2</type>
<position>40,-85.5</position>
<input>
<ID>IN_0</ID>216 </input>
<input>
<ID>IN_1</ID>217 </input>
<output>
<ID>OUT</ID>219 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>376</ID>
<type>BA_NAND2</type>
<position>41.5,-98.5</position>
<input>
<ID>IN_0</ID>216 </input>
<input>
<ID>IN_1</ID>215 </input>
<output>
<ID>OUT</ID>221 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>378</ID>
<type>BA_NAND2</type>
<position>49.5,-79</position>
<input>
<ID>IN_0</ID>218 </input>
<input>
<ID>IN_1</ID>219 </input>
<output>
<ID>OUT</ID>220 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>380</ID>
<type>GA_LED</type>
<position>60,-79</position>
<input>
<ID>N_in0</ID>220 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>381</ID>
<type>GA_LED</type>
<position>49,-99.5</position>
<input>
<ID>N_in0</ID>221 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>383</ID>
<type>AA_LABEL</type>
<position>69,-87.5</position>
<gparam>LABEL_TEXT redesign</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>202</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-35,28.5,-1</points>
<intersection>-35 3</intersection>
<intersection>-8 2</intersection>
<intersection>-1 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,-1,40,-1</points>
<connection>
<GID>351</GID>
<name>IN_0</name></connection>
<intersection>28.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-8,28.5,-8</points>
<connection>
<GID>347</GID>
<name>OUT_0</name></connection>
<intersection>28.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>28.5,-35,40,-35</points>
<connection>
<GID>353</GID>
<name>IN_0</name></connection>
<intersection>28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,-27,15,-3</points>
<intersection>-27 1</intersection>
<intersection>-27 1</intersection>
<intersection>-3 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6.5,-27,19,-27</points>
<connection>
<GID>348</GID>
<name>IN_0</name></connection>
<connection>
<GID>358</GID>
<name>OUT_0</name></connection>
<intersection>15 0</intersection>
<intersection>16.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15,-3,40,-3</points>
<connection>
<GID>351</GID>
<name>IN_1</name></connection>
<intersection>15 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>16.5,-37,16.5,-27</points>
<intersection>-37 4</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>16.5,-37,40,-37</points>
<connection>
<GID>353</GID>
<name>IN_1</name></connection>
<intersection>16.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-16.5,18,-8</points>
<intersection>-16.5 2</intersection>
<intersection>-9.5 3</intersection>
<intersection>-8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-8,19,-8</points>
<connection>
<GID>347</GID>
<name>IN_0</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18,-16.5,40.5,-16.5</points>
<connection>
<GID>352</GID>
<name>IN_0</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>5.5,-9.5,18,-9.5</points>
<connection>
<GID>357</GID>
<name>OUT_0</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-27,32.5,-18.5</points>
<intersection>-27 1</intersection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-27,32.5,-27</points>
<connection>
<GID>348</GID>
<name>OUT_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-18.5,40.5,-18.5</points>
<connection>
<GID>352</GID>
<name>IN_1</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-8.5,50.5,-2</points>
<intersection>-8.5 1</intersection>
<intersection>-2 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-8.5,55,-8.5</points>
<connection>
<GID>355</GID>
<name>IN_0</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46,-2,50.5,-2</points>
<connection>
<GID>351</GID>
<name>OUT</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-17.5,50.5,-10.5</points>
<intersection>-17.5 2</intersection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-10.5,55,-10.5</points>
<connection>
<GID>355</GID>
<name>IN_1</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46.5,-17.5,50.5,-17.5</points>
<connection>
<GID>352</GID>
<name>OUT</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61,-9.5,63.5,-9.5</points>
<connection>
<GID>360</GID>
<name>N_in0</name></connection>
<connection>
<GID>355</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>209</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-36.5,47,-36</points>
<intersection>-36.5 1</intersection>
<intersection>-36 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-36.5,48,-36.5</points>
<connection>
<GID>361</GID>
<name>N_in0</name></connection>
<intersection>47 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46,-36,47,-36</points>
<connection>
<GID>353</GID>
<name>OUT</name></connection>
<intersection>47 0</intersection></hsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,-94.5,6,-70</points>
<intersection>-94.5 3</intersection>
<intersection>-94 1</intersection>
<intersection>-92.5 4</intersection>
<intersection>-70 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1,-94,6,-94</points>
<connection>
<GID>365</GID>
<name>OUT_0</name></connection>
<intersection>6 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>6,-70,35.5,-70</points>
<intersection>6 0</intersection>
<intersection>35.5 5</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>6,-94.5,14,-94.5</points>
<connection>
<GID>372</GID>
<name>IN_1</name></connection>
<intersection>6 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>6,-92.5,14,-92.5</points>
<connection>
<GID>372</GID>
<name>IN_0</name></connection>
<intersection>6 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>35.5,-99.5,35.5,-70</points>
<intersection>-99.5 7</intersection>
<intersection>-75.5 8</intersection>
<intersection>-70 2</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>35.5,-99.5,38.5,-99.5</points>
<connection>
<GID>376</GID>
<name>IN_1</name></connection>
<intersection>35.5 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>35.5,-75.5,38.5,-75.5</points>
<connection>
<GID>374</GID>
<name>IN_1</name></connection>
<intersection>35.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>216</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-97.5,30,-73.5</points>
<intersection>-97.5 3</intersection>
<intersection>-84.5 4</intersection>
<intersection>-75.5 2</intersection>
<intersection>-73.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-73.5,38.5,-73.5</points>
<connection>
<GID>374</GID>
<name>IN_0</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21.5,-75.5,30,-75.5</points>
<connection>
<GID>371</GID>
<name>OUT</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>30,-97.5,38.5,-97.5</points>
<connection>
<GID>376</GID>
<name>IN_0</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>30,-84.5,37,-84.5</points>
<connection>
<GID>375</GID>
<name>IN_0</name></connection>
<intersection>30 0</intersection></hsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-93.5,28.5,-86.5</points>
<intersection>-93.5 1</intersection>
<intersection>-86.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20,-93.5,28.5,-93.5</points>
<connection>
<GID>372</GID>
<name>OUT</name></connection>
<intersection>28.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-86.5,37,-86.5</points>
<connection>
<GID>375</GID>
<name>IN_1</name></connection>
<intersection>28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,-78,45.5,-74.5</points>
<intersection>-78 1</intersection>
<intersection>-74.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45.5,-78,46.5,-78</points>
<connection>
<GID>378</GID>
<name>IN_0</name></connection>
<intersection>45.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>44.5,-74.5,45.5,-74.5</points>
<connection>
<GID>374</GID>
<name>OUT</name></connection>
<intersection>45.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-85.5,44.5,-80</points>
<intersection>-85.5 2</intersection>
<intersection>-80 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44.5,-80,46.5,-80</points>
<connection>
<GID>378</GID>
<name>IN_1</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43,-85.5,44.5,-85.5</points>
<connection>
<GID>375</GID>
<name>OUT</name></connection>
<intersection>44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>52.5,-79,59,-79</points>
<connection>
<GID>380</GID>
<name>N_in0</name></connection>
<connection>
<GID>378</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-99.5,46,-98.5</points>
<intersection>-99.5 1</intersection>
<intersection>-98.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-99.5,48,-99.5</points>
<connection>
<GID>381</GID>
<name>N_in0</name></connection>
<intersection>46 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>44.5,-98.5,46,-98.5</points>
<connection>
<GID>376</GID>
<name>OUT</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15.5,-76.5,15.5,-74.5</points>
<connection>
<GID>371</GID>
<name>IN_1</name></connection>
<connection>
<GID>371</GID>
<name>IN_0</name></connection>
<intersection>-75.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1,-75.5,15.5,-75.5</points>
<connection>
<GID>364</GID>
<name>OUT_0</name></connection>
<intersection>15.5 0</intersection></hsegment></shape></wire></page 5>
<page 6>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 9></circuit>